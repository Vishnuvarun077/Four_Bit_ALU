magic
tech scmos
timestamp 1700591413
<< nwell >>
rect 180 59 270 77
rect 416 70 506 88
rect 305 -56 342 -38
rect 348 -56 372 -38
rect 433 -55 470 -37
rect 476 -55 500 -37
rect 474 -127 531 -109
<< ntransistor >>
rect 191 19 193 23
rect 207 19 209 23
rect 217 19 219 23
rect 227 19 229 23
rect 237 19 239 23
rect 427 30 429 34
rect 443 30 445 34
rect 453 30 455 34
rect 463 30 465 34
rect 473 30 475 34
rect 257 19 259 23
rect 493 30 495 34
rect 316 -80 318 -76
rect 326 -80 328 -76
rect 359 -80 361 -76
rect 444 -79 446 -75
rect 454 -79 456 -75
rect 487 -79 489 -75
rect 485 -157 487 -153
rect 495 -157 497 -153
rect 513 -157 515 -153
<< ptransistor >>
rect 191 65 193 71
rect 207 65 209 71
rect 217 65 219 71
rect 227 65 229 71
rect 237 65 239 71
rect 257 65 259 71
rect 427 76 429 82
rect 443 76 445 82
rect 453 76 455 82
rect 463 76 465 82
rect 473 76 475 82
rect 493 76 495 82
rect 316 -50 318 -44
rect 326 -50 328 -44
rect 359 -50 361 -44
rect 444 -49 446 -43
rect 454 -49 456 -43
rect 487 -49 489 -43
rect 485 -121 487 -115
rect 495 -121 497 -115
rect 513 -121 515 -115
<< ndiffusion >>
rect 190 19 191 23
rect 193 19 194 23
rect 206 19 207 23
rect 209 19 217 23
rect 219 19 221 23
rect 225 19 227 23
rect 229 19 237 23
rect 239 19 240 23
rect 426 30 427 34
rect 429 30 430 34
rect 442 30 443 34
rect 445 30 453 34
rect 455 30 457 34
rect 461 30 463 34
rect 465 30 473 34
rect 475 30 476 34
rect 256 19 257 23
rect 259 19 260 23
rect 492 30 493 34
rect 495 30 496 34
rect 315 -80 316 -76
rect 318 -80 326 -76
rect 328 -80 330 -76
rect 358 -80 359 -76
rect 361 -80 362 -76
rect 443 -79 444 -75
rect 446 -79 454 -75
rect 456 -79 458 -75
rect 486 -79 487 -75
rect 489 -79 490 -75
rect 484 -157 485 -153
rect 487 -157 489 -153
rect 493 -157 495 -153
rect 497 -157 498 -153
rect 512 -157 513 -153
rect 515 -157 516 -153
<< pdiffusion >>
rect 190 65 191 71
rect 193 65 194 71
rect 206 65 207 71
rect 209 65 217 71
rect 219 65 221 71
rect 225 65 227 71
rect 229 65 237 71
rect 239 65 240 71
rect 256 65 257 71
rect 259 65 260 71
rect 426 76 427 82
rect 429 76 430 82
rect 442 76 443 82
rect 445 76 453 82
rect 455 76 457 82
rect 461 76 463 82
rect 465 76 473 82
rect 475 76 476 82
rect 492 76 493 82
rect 495 76 496 82
rect 315 -50 316 -44
rect 318 -50 320 -44
rect 324 -50 326 -44
rect 328 -50 330 -44
rect 358 -50 359 -44
rect 361 -50 362 -44
rect 443 -49 444 -43
rect 446 -49 448 -43
rect 452 -49 454 -43
rect 456 -49 458 -43
rect 486 -49 487 -43
rect 489 -49 490 -43
rect 484 -121 485 -115
rect 487 -121 495 -115
rect 497 -121 498 -115
rect 512 -121 513 -115
rect 515 -121 516 -115
<< ndcontact >>
rect 186 19 190 23
rect 194 19 198 23
rect 202 19 206 23
rect 221 19 225 23
rect 240 19 244 23
rect 422 30 426 34
rect 430 30 434 34
rect 438 30 442 34
rect 457 30 461 34
rect 476 30 480 34
rect 252 19 256 23
rect 260 19 264 23
rect 488 30 492 34
rect 496 30 500 34
rect 311 -80 315 -76
rect 330 -80 334 -76
rect 354 -80 358 -76
rect 362 -80 366 -76
rect 439 -79 443 -75
rect 458 -79 462 -75
rect 482 -79 486 -75
rect 490 -79 494 -75
rect 480 -157 484 -153
rect 489 -157 493 -153
rect 498 -157 502 -153
rect 508 -157 512 -153
rect 516 -157 520 -153
<< pdcontact >>
rect 186 65 190 71
rect 194 65 198 71
rect 202 65 206 71
rect 221 65 225 71
rect 240 65 244 71
rect 252 65 256 71
rect 260 65 264 71
rect 422 76 426 82
rect 430 76 434 82
rect 438 76 442 82
rect 457 76 461 82
rect 476 76 480 82
rect 488 76 492 82
rect 496 76 500 82
rect 311 -50 315 -44
rect 320 -50 324 -44
rect 330 -50 334 -44
rect 354 -50 358 -44
rect 362 -50 366 -44
rect 439 -49 443 -43
rect 448 -49 452 -43
rect 458 -49 462 -43
rect 482 -49 486 -43
rect 490 -49 494 -43
rect 480 -121 484 -115
rect 498 -121 502 -115
rect 508 -121 512 -115
rect 516 -121 520 -115
<< polysilicon >>
rect 427 90 513 92
rect 427 82 429 90
rect 443 82 445 85
rect 453 82 455 85
rect 463 82 465 90
rect 473 82 475 85
rect 493 82 495 85
rect 191 79 277 81
rect 191 71 193 79
rect 207 71 209 74
rect 217 71 219 74
rect 227 71 229 79
rect 237 71 239 74
rect 257 71 259 74
rect 191 23 193 65
rect 207 23 209 65
rect 217 44 219 65
rect 227 62 229 65
rect 217 42 229 44
rect 217 23 219 26
rect 227 23 229 42
rect 237 23 239 65
rect 257 42 259 65
rect 275 37 277 79
rect 248 35 277 37
rect 191 16 193 19
rect 207 8 209 19
rect 217 13 219 19
rect 227 16 229 19
rect 237 16 239 19
rect 248 13 250 35
rect 427 34 429 76
rect 443 34 445 76
rect 453 55 455 76
rect 463 73 465 76
rect 453 53 465 55
rect 453 34 455 37
rect 463 34 465 53
rect 473 34 475 76
rect 493 53 495 76
rect 511 48 513 90
rect 484 46 513 48
rect 257 23 259 31
rect 427 27 429 30
rect 443 19 445 30
rect 453 24 455 30
rect 463 27 465 30
rect 473 27 475 30
rect 484 24 486 46
rect 493 34 495 42
rect 453 22 486 24
rect 493 19 495 30
rect 217 11 250 13
rect 257 8 259 19
rect 443 17 495 19
rect 207 6 259 8
rect 316 -44 318 -35
rect 326 -44 328 -35
rect 359 -44 361 -35
rect 444 -43 446 -34
rect 454 -43 456 -34
rect 487 -43 489 -34
rect 316 -76 318 -50
rect 326 -76 328 -50
rect 359 -76 361 -50
rect 444 -75 446 -49
rect 454 -75 456 -49
rect 487 -75 489 -49
rect 316 -83 318 -80
rect 326 -83 328 -80
rect 359 -83 361 -80
rect 444 -82 446 -79
rect 454 -82 456 -79
rect 487 -82 489 -79
rect 485 -115 487 -112
rect 495 -115 497 -112
rect 513 -115 515 -112
rect 485 -153 487 -121
rect 495 -153 497 -121
rect 513 -153 515 -121
rect 485 -160 487 -157
rect 495 -160 497 -157
rect 513 -160 515 -157
<< polycontact >>
rect 187 42 191 46
rect 213 42 217 46
rect 239 42 243 46
rect 259 42 263 46
rect 423 53 427 57
rect 449 53 453 57
rect 475 53 479 57
rect 495 53 499 57
rect 259 27 263 31
rect 495 38 499 42
rect 312 -62 316 -58
rect 322 -71 326 -67
rect 355 -62 359 -58
rect 440 -61 444 -57
rect 450 -70 454 -66
rect 483 -61 487 -57
rect 481 -134 485 -130
rect 491 -141 495 -137
rect 509 -139 513 -135
<< metal1 >>
rect 387 95 553 99
rect 387 90 392 95
rect 300 89 392 90
rect 266 88 392 89
rect 180 85 392 88
rect 180 84 306 85
rect 186 71 190 84
rect 202 71 206 84
rect 240 71 244 84
rect 260 71 264 84
rect 422 82 426 95
rect 438 82 442 95
rect 476 82 480 95
rect 496 82 500 95
rect 547 94 553 95
rect 129 46 185 47
rect 194 46 198 65
rect 221 55 225 65
rect 129 42 187 46
rect 194 42 213 46
rect 129 33 137 39
rect 129 -9 144 -3
rect 154 -58 160 42
rect 194 23 198 42
rect 221 23 225 50
rect 252 46 256 65
rect 300 54 399 57
rect 287 53 399 54
rect 430 57 434 76
rect 457 66 461 76
rect 404 53 423 57
rect 430 53 449 57
rect 287 50 304 53
rect 243 42 256 46
rect 252 23 256 42
rect 263 39 267 46
rect 263 27 267 34
rect 392 45 416 49
rect 186 5 190 19
rect 202 5 206 19
rect 240 5 244 19
rect 260 5 264 19
rect 300 5 306 7
rect 181 1 306 5
rect 276 -4 281 -3
rect 392 -4 396 45
rect 430 34 434 53
rect 457 34 461 61
rect 488 57 492 76
rect 569 61 575 66
rect 479 53 492 57
rect 488 34 492 53
rect 499 50 503 57
rect 499 38 503 45
rect 422 17 426 30
rect 417 16 426 17
rect 438 16 442 30
rect 476 16 480 30
rect 496 16 500 30
rect 417 12 507 16
rect 180 -8 396 -4
rect 369 -26 374 -24
rect 305 -29 374 -26
rect 311 -44 315 -29
rect 330 -44 334 -29
rect 354 -44 358 -29
rect 320 -58 324 -50
rect 362 -58 366 -50
rect 392 -57 396 -8
rect 428 -25 433 -24
rect 524 -25 532 -24
rect 428 -28 554 -25
rect 428 -29 433 -28
rect 439 -43 443 -28
rect 458 -43 462 -28
rect 482 -43 486 -28
rect 524 -29 532 -28
rect 448 -57 452 -49
rect 490 -57 494 -49
rect 372 -58 385 -57
rect 154 -62 312 -58
rect 320 -62 355 -58
rect 362 -62 385 -58
rect 392 -61 440 -57
rect 448 -61 483 -57
rect 490 -61 547 -57
rect 155 -63 304 -62
rect 284 -71 322 -67
rect 330 -76 334 -62
rect 362 -76 366 -62
rect 276 -86 281 -85
rect 276 -87 306 -86
rect 311 -87 315 -80
rect 354 -87 358 -80
rect 368 -87 373 -85
rect 276 -90 373 -87
rect 378 -137 385 -62
rect 404 -70 450 -66
rect 458 -75 462 -61
rect 490 -75 494 -61
rect 431 -86 436 -85
rect 439 -86 443 -79
rect 482 -86 486 -79
rect 431 -89 501 -86
rect 431 -90 436 -89
rect 474 -103 532 -98
rect 480 -115 484 -103
rect 508 -115 512 -103
rect 524 -104 532 -103
rect 434 -134 481 -130
rect 434 -178 438 -134
rect 498 -135 502 -121
rect 516 -135 520 -121
rect 477 -141 491 -137
rect 498 -139 509 -135
rect 516 -139 532 -135
rect 498 -145 502 -139
rect 489 -149 502 -145
rect 489 -153 493 -149
rect 516 -153 520 -139
rect 480 -164 484 -157
rect 498 -164 502 -157
rect 508 -164 512 -157
rect 467 -169 530 -164
rect 543 -178 547 -61
rect 571 -139 576 -134
rect 434 -183 547 -178
<< m2contact >>
rect 221 50 226 55
rect 137 33 144 39
rect 282 50 287 55
rect 399 53 404 58
rect 457 61 462 66
rect 262 34 267 39
rect 416 45 421 50
rect 564 61 569 66
rect 498 45 503 50
rect 276 -73 284 -66
rect 399 -70 404 -65
rect 378 -143 386 -137
rect 470 -143 477 -137
rect 532 -139 537 -134
rect 566 -139 571 -134
<< metal2 >>
rect 462 61 564 65
rect 226 50 282 54
rect 144 34 262 39
rect 144 33 172 34
rect 166 -66 172 33
rect 399 -65 404 53
rect 421 45 498 50
rect 166 -73 276 -66
rect 399 -71 404 -70
rect 386 -143 470 -137
rect 537 -139 566 -135
<< m3contact >>
rect 547 94 553 99
rect 136 -9 144 -3
rect 300 1 306 7
rect 180 -9 185 -3
rect 276 -8 281 -3
rect 369 -29 374 -24
rect 417 12 422 17
rect 428 -29 433 -24
rect 524 -29 532 -24
rect 547 -28 554 -23
rect 276 -90 281 -85
rect 368 -90 373 -85
rect 431 -90 436 -85
rect 524 -104 532 -98
rect 466 -169 472 -164
<< metal3 >>
rect 417 7 422 12
rect 306 3 422 7
rect 276 -3 281 -2
rect 144 -9 180 -3
rect 276 -85 281 -8
rect 547 -23 553 94
rect 374 -29 428 -25
rect 433 -29 436 -25
rect 373 -90 431 -87
rect 404 -164 408 -90
rect 524 -98 531 -29
rect 404 -169 466 -164
rect 472 -169 476 -164
<< labels >>
rlabel metal1 305 -29 372 -26 1 VDD
rlabel metal1 304 -90 373 -87 1 GND
rlabel metal1 470 -134 478 -130 1 t2
rlabel metal1 470 -141 478 -137 1 t1
rlabel metal1 569 61 575 66 7 SUM
rlabel metal1 571 -139 576 -134 7 COUT
rlabel metal1 129 42 135 47 3 B
rlabel metal1 129 33 137 39 3 A
rlabel metal1 129 -9 136 -3 3 Cin
rlabel metal1 204 84 209 88 1 VDD
rlabel metal1 270 1 275 5 1 GND
rlabel metal1 287 -71 292 -67 1 A
rlabel metal1 284 -63 289 -59 1 B
rlabel metal1 472 95 477 99 5 VDD
rlabel metal1 460 12 465 16 1 GND
rlabel metal1 391 -8 396 -4 1 Cin
rlabel metal1 390 53 395 57 1 D1
rlabel metal1 449 -28 455 -25 1 VDD
rlabel metal1 455 -89 461 -86 1 GND
rlabel metal1 494 -101 500 -98 1 VDD
rlabel metal1 491 -168 497 -165 1 GND
<< end >>
