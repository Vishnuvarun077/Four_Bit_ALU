magic
tech scmos
timestamp 1699212410
<< nwell >>
rect -25 -4 65 14
<< polysilicon >>
rect -14 16 72 18
rect -14 8 -12 16
rect 2 8 4 11
rect 12 8 14 11
rect 22 8 24 16
rect 32 8 34 11
rect 52 8 54 11
rect -14 -40 -12 2
rect 2 -40 4 2
rect 12 -19 14 2
rect 22 -1 24 2
rect 12 -21 24 -19
rect 12 -40 14 -37
rect 22 -40 24 -21
rect 32 -40 34 2
rect 52 -21 54 2
rect 70 -26 72 16
rect 43 -28 72 -26
rect -14 -47 -12 -44
rect 2 -55 4 -44
rect 12 -50 14 -44
rect 22 -47 24 -44
rect 32 -47 34 -44
rect 43 -50 45 -28
rect 52 -40 54 -32
rect 12 -52 45 -50
rect 52 -55 54 -44
rect 2 -57 54 -55
<< ndiffusion >>
rect -15 -44 -14 -40
rect -12 -44 -11 -40
rect 1 -44 2 -40
rect 4 -44 12 -40
rect 14 -44 16 -40
rect 20 -44 22 -40
rect 24 -44 32 -40
rect 34 -44 35 -40
rect 51 -44 52 -40
rect 54 -44 55 -40
<< pdiffusion >>
rect -15 2 -14 8
rect -12 2 -11 8
rect 1 2 2 8
rect 4 2 12 8
rect 14 2 16 8
rect 20 2 22 8
rect 24 2 32 8
rect 34 2 35 8
rect 51 2 52 8
rect 54 2 55 8
<< metal1 >>
rect -25 21 65 25
rect -19 8 -15 21
rect -3 8 1 21
rect 35 8 39 21
rect 55 8 59 21
rect -11 -17 -7 2
rect 16 -8 20 2
rect -33 -21 -18 -17
rect -11 -21 8 -17
rect -33 -29 -25 -25
rect -11 -40 -7 -21
rect 16 -40 20 -13
rect 47 -17 51 2
rect 82 -13 91 -9
rect 38 -21 51 -17
rect 47 -40 51 -21
rect 58 -24 62 -17
rect 58 -36 62 -29
rect -19 -58 -15 -44
rect -3 -58 1 -44
rect 35 -58 39 -44
rect 55 -58 59 -44
rect -24 -62 66 -58
<< metal2 >>
rect 21 -13 77 -9
rect -20 -29 57 -24
<< ntransistor >>
rect -14 -44 -12 -40
rect 2 -44 4 -40
rect 12 -44 14 -40
rect 22 -44 24 -40
rect 32 -44 34 -40
rect 52 -44 54 -40
<< ptransistor >>
rect -14 2 -12 8
rect 2 2 4 8
rect 12 2 14 8
rect 22 2 24 8
rect 32 2 34 8
rect 52 2 54 8
<< polycontact >>
rect -18 -21 -14 -17
rect 8 -21 12 -17
rect 34 -21 38 -17
rect 54 -21 58 -17
rect 54 -36 58 -32
<< ndcontact >>
rect -19 -44 -15 -40
rect -11 -44 -7 -40
rect -3 -44 1 -40
rect 16 -44 20 -40
rect 35 -44 39 -40
rect 47 -44 51 -40
rect 55 -44 59 -40
<< pdcontact >>
rect -19 2 -15 8
rect -11 2 -7 8
rect -3 2 1 8
rect 16 2 20 8
rect 35 2 39 8
rect 47 2 51 8
rect 55 2 59 8
<< m2contact >>
rect 16 -13 21 -8
rect -25 -29 -20 -24
rect 77 -13 82 -8
rect 57 -29 62 -24
<< labels >>
rlabel metal1 -25 21 65 25 5 VDD
rlabel metal1 -33 -21 -14 -17 1 B
rlabel metal1 -11 -21 12 -17 1 Bnot
rlabel metal1 -24 -62 66 -58 1 GND
rlabel space -33 -29 62 -25 1 A
rlabel metal1 34 -21 46 -17 1 Anot
rlabel metal2 16 -13 82 -9 1 XOR
rlabel metal1 16 -44 20 8 1 xor
rlabel metal1 16 -44 20 8 1 XOR
rlabel metal1 54 -21 62 -17 1 A
rlabel metal1 54 -36 62 -32 1 A
<< end >>
