magic
tech scmos
timestamp 1699022636
<< nwell >>
rect -9 1 16 17
<< polysilicon >>
rect 2 11 4 14
rect 2 -2 4 7
rect -2 -4 4 -2
rect 2 -9 4 -4
rect 2 -16 4 -13
<< ndiffusion >>
rect 1 -13 2 -9
rect 4 -13 5 -9
<< pdiffusion >>
rect 1 7 2 11
rect 4 7 5 11
<< metal1 >>
rect -9 17 16 20
rect -2 11 1 17
rect -8 -5 -6 -1
rect 5 -2 8 7
rect 5 -5 16 -2
rect 5 -9 8 -5
rect -2 -17 1 -13
rect -9 -20 16 -17
<< ntransistor >>
rect 2 -13 4 -9
<< ptransistor >>
rect 2 7 4 11
<< polycontact >>
rect -6 -5 -2 -1
<< ndcontact >>
rect -3 -13 1 -9
rect 5 -13 9 -9
<< pdcontact >>
rect -3 7 1 11
rect 5 7 9 11
<< labels >>
rlabel metal1 -2 -19 0 -18 1 gnd
rlabel metal1 -5 18 -3 19 4 vdd
rlabel metal1 -8 -4 -7 -2 3 input
rlabel metal1 14 -4 16 -3 7 output
<< end >>
