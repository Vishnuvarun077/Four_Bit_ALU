* SPICE3 file created from comparatorfinal.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8V
.option scale=0.09u
Vds VDD GND 'SUPPLY'


* V_in_a3 CompA3 GND PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
* V_in_a2 CompA2 GND PULSE(0 1.8 0ns 100ps 100ps 30ns 50ns)
* V_in_a1 CompA1 GND PULSE(0 1.8 0ns 100ps 100ps 40ns 60ns)
* V_in_a0 CompA0 GND PULSE(0 1.8 0ns 100ps 100ps 50ns 80ns)

*  V_in_b3 CompB3 GND PULSE(0 1.8 0ns 100ps 100ps 10ns 50ns)
*  V_in_b2 CompB2 GND PULSE(0 1.8 0ns 100ps 100ps 20ns 60ns)
* V_in_b1 CompB1 GND PULSE(0 1.8 0ns 100ps 100ps 30ns 70ns)
* V_in_b0 CompB0 GND PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
V_in_a3 CompA3 GND PULSE(0 1.8 0ns 100ps 100ps 10ns 40ns)
V_in_a2 CompA2 GND PULSE(0 1.8 0ns 100ps 100ps 20ns 50ns)
V_in_a1 CompA1 GND PULSE(0 1.8 0ns 100ps 100ps 30ns 60ns)
V_in_a0 CompA0 GND PULSE(0 1.8 0ns 100ps 100ps 40ns 70ns)

V_in_b3 CompB3 GND PULSE(0 1.8 0ns 100ps 100ps 50ns 90ns)
V_in_b2 CompB2 GND PULSE(0 1.8 0ns 100ps 100ps 60ns 100ns)
V_in_b1 CompB1 GND PULSE(0 1.8 0ns 100ps 100ps 70ns 110ns)
V_in_b0 CompB0 GND PULSE(0 1.8 0ns 100ps 100ps 80ns 120ns)


.option scale=0.09u

M1000 VDD n2 a_16444_n18992# w_16431_n18998# CMOSP w=6 l=2
+  ad=1378 pd=994 as=96 ps=56
M1001 a_15971_n19304# CompA1 a_15991_n19345# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1002 AGB a_16493_n19415# VDD w_16480_n19371# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1003 a_16262_n19342# CompA0 a_16252_n19342# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1004 a_16444_n18992# n3 VDD w_16431_n18998# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_15991_n19345# CompB1not a_15981_n19345# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1006 a_15449_n19164# CompA3 VDD w_15436_n19124# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1007 a_16252_n19342# n1 a_16242_n19342# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1008 a_15449_n19164# CompA3 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=812 ps=726
M1009 a_15981_n19345# n2 a_15971_n19345# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1010 VDD CompB2 a_15742_n19167# w_15685_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=30 ps=22
M1011 a_16242_n19342# n2 a_16232_n19342# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1012 a_15514_n19318# CompB3not a_15514_n19348# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1013 y2 a_15716_n19313# VDD w_15756_n19319# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1014 GND CompB2 a_15742_n19167# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1015 CompB3not CompB3 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1016 a_15971_n19345# n3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 y0 a_16232_n19294# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1018 a_16232_n19342# n3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 a_15514_n19348# CompA3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 VDD a_15742_n19167# a_15734_n19118# w_15685_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1021 CompB0not CompB0 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1022 GND a_15742_n19167# a_15734_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1023 a_15734_n19118# CompA2 a_15724_n19164# w_15685_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1024 CompB2not CompB2 VDD w_15617_n19485# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1025 a_15734_n19164# a_15698_n19164# a_15724_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1026 a_15724_n19164# a_15698_n19164# a_15714_n19118# w_15685_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1027 a_15724_n19164# CompA2 a_15714_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1028 a_15714_n19118# CompB2 VDD w_15685_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 a_16177_n19164# CompA0 VDD w_16164_n19124# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1030 a_15714_n19164# CompB2 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 a_16177_n19164# CompA0 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1032 ALB AGB a_16743_n19147# w_16730_n19153# CMOSP w=6 l=2
+  ad=30 pd=22 as=48 ps=28
M1033 a_16743_n19147# AEB VDD w_16730_n19153# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 VDD CompA1 a_15971_n19304# w_15958_n19310# CMOSP w=6 l=2
+  ad=0 pd=0 as=96 ps=56
M1035 AEB a_16444_n18992# VDD w_16492_n18998# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1036 a_16493_n19415# y3 GND Gnd CMOSN w=4 l=2
+  ad=64 pd=48 as=0 ps=0
M1037 a_15971_n19304# CompB1not VDD w_15958_n19310# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 n0 a_16203_n19164# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1039 VDD n2 a_15971_n19304# w_15958_n19310# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 VDD a_15493_n19167# a_15485_n19118# w_15436_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1041 a_15971_n19304# n3 VDD w_15958_n19310# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 GND a_15493_n19167# a_15485_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1043 a_15485_n19118# CompA3 a_15475_n19164# w_15436_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1044 a_15485_n19164# a_15449_n19164# a_15475_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1045 a_16444_n18992# n0 a_16464_n19033# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1046 y3 a_15514_n19318# VDD w_15544_n19324# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1047 a_15475_n19164# a_15449_n19164# a_15465_n19118# w_15436_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1048 a_15475_n19164# CompA3 a_15465_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1049 a_16464_n19033# n1 a_16454_n19033# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1050 a_15465_n19118# CompB3 VDD w_15436_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 a_15465_n19164# CompB3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 CompB3not CompB3 VDD w_15561_n19485# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1053 a_16454_n19033# n2 a_16444_n19033# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1054 a_16444_n19033# n3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 a_15955_n19164# CompA1 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1056 a_15955_n19164# CompA1 VDD w_15942_n19124# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1057 CompB0not CompB0 VDD w_16077_n19485# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1058 a_16493_n19365# y3 VDD w_16480_n19371# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1059 a_15716_n19313# CompA2 VDD w_15703_n19319# CMOSP w=6 l=2
+  ad=84 pd=52 as=0 ps=0
M1060 a_15698_n19164# CompA2 VDD w_15685_n19124# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1061 VDD CompB2not a_15716_n19313# w_15703_n19319# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 a_15698_n19164# CompA2 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1063 a_15716_n19313# n3 VDD w_15703_n19319# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 a_16193_n19118# CompB0 VDD w_16164_n19124# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1065 GND AGB ALB Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1066 a_16193_n19164# CompB0 GND Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1067 n2 a_15724_n19164# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1068 CompB1not CompB1 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1069 ALB AEB GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 y2 a_15716_n19313# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1071 a_16232_n19294# CompB0not VDD w_16219_n19300# CMOSP w=6 l=2
+  ad=132 pd=80 as=0 ps=0
M1072 n0 a_16203_n19164# VDD w_16304_n19127# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1073 VDD CompA0 a_16232_n19294# w_16219_n19300# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 AEB a_16444_n18992# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1075 a_16232_n19294# n1 VDD w_16219_n19300# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 VDD n2 a_16232_n19294# w_16219_n19300# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 GND y2 a_16493_n19415# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 y0 a_16232_n19294# VDD w_16292_n19300# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1079 a_16232_n19294# n3 VDD w_16219_n19300# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 n1 a_15981_n19164# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1081 VDD CompB3 a_15493_n19167# w_15436_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=30 ps=22
M1082 VDD CompB3not a_15514_n19318# w_15501_n19324# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1083 GND CompB3 a_15493_n19167# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1084 GND y0 a_16493_n19415# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 n3 a_15475_n19164# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1086 a_15514_n19318# CompA3 VDD w_15501_n19324# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 a_16493_n19415# y1 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 y3 a_15514_n19318# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1089 GND CompB1 a_15999_n19167# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1090 VDD CompB1 a_15999_n19167# w_15942_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=30 ps=22
M1091 y1 a_15971_n19304# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1092 VDD a_15999_n19167# a_15991_n19118# w_15942_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1093 GND a_15999_n19167# a_15991_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1094 a_15991_n19118# CompA1 a_15981_n19164# w_15942_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1095 a_15991_n19164# a_15955_n19164# a_15981_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1096 VDD CompB0 a_16221_n19167# w_16164_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=30 ps=22
M1097 a_15981_n19164# a_15955_n19164# a_15971_n19118# w_15942_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1098 n2 a_15724_n19164# VDD w_15825_n19127# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1099 CompB1not CompB1 VDD w_15814_n19485# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1100 a_16503_n19365# y2 a_16493_n19365# w_16480_n19371# CMOSP w=6 l=2
+  ad=42 pd=26 as=0 ps=0
M1101 GND CompB0 a_16221_n19167# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1102 a_15981_n19164# CompA1 a_15971_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1103 a_15971_n19118# CompB1 VDD w_15942_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 CompB2not CompB2 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1105 a_15971_n19164# CompB1 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 AGB a_16493_n19415# GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1107 VDD a_16221_n19167# a_16213_n19118# w_16164_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1108 a_16493_n19415# y0 a_16512_n19365# w_16480_n19371# CMOSP w=6 l=2
+  ad=36 pd=24 as=48 ps=28
M1109 GND a_16221_n19167# a_16213_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1110 a_16213_n19118# CompA0 a_16203_n19164# w_16164_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1111 a_16512_n19365# y1 a_16503_n19365# w_16480_n19371# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 a_15716_n19313# CompA2 a_15726_n19346# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1113 a_16213_n19164# a_16177_n19164# a_16203_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1114 a_16203_n19164# CompA0 a_16193_n19164# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 a_16203_n19164# a_16177_n19164# a_16193_n19118# w_16164_n19124# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 a_15726_n19346# CompB2not a_15716_n19346# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1117 a_15716_n19346# n3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 n1 a_15981_n19164# VDD w_16082_n19127# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1119 VDD n0 a_16444_n18992# w_16431_n18998# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 y1 a_15971_n19304# VDD w_16019_n19310# CMOSP w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1121 a_16444_n18992# n1 VDD w_16431_n18998# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 n3 a_15475_n19164# VDD w_15576_n19127# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1123 a_16232_n19294# CompB0not a_16262_n19342# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
C0 GND VDD 0.43fF
C1 CompB3not w_15561_n19485# 0.03fF
C2 VDD n1 0.38fF
C3 a_15955_n19164# GND 0.08fF
C4 y1 VDD 0.06fF
C5 CompA0 w_16164_n19124# 0.14fF
C6 w_16304_n19127# n0 0.03fF
C7 a_16203_n19164# w_16304_n19127# 0.06fF
C8 n2 w_15958_n19310# 0.08fF
C9 a_15716_n19313# VDD 0.13fF
C10 n3 a_15475_n19164# 0.02fF
C11 AEB w_16492_n18998# 0.03fF
C12 w_15703_n19319# VDD 0.05fF
C13 a_16203_n19164# w_16164_n19124# 0.02fF
C14 w_15825_n19127# VDD 0.05fF
C15 CompB3not CompB3 0.02fF
C16 CompB0not y3 0.10fF
C17 w_15685_n19124# CompB2 0.13fF
C18 w_15544_n19324# VDD 0.03fF
C19 CompA0 n3 0.18fF
C20 w_15685_n19124# VDD 0.12fF
C21 GND n2 0.17fF
C22 a_15698_n19164# CompA2 0.08fF
C23 n3 w_15576_n19127# 0.03fF
C24 n3 n0 0.08fF
C25 n2 n1 6.42fF
C26 a_15724_n19164# CompA2 0.01fF
C27 y3 y2 9.36fF
C28 CompB0not CompA0 0.57fF
C29 GND a_16232_n19294# 0.02fF
C30 w_16077_n19485# VDD 0.05fF
C31 VDD CompB2 0.24fF
C32 CompB1not VDD 0.15fF
C33 a_16232_n19294# n1 0.08fF
C34 CompB1not w_15814_n19485# 0.03fF
C35 w_15814_n19485# VDD 0.05fF
C36 AGB a_16493_n19415# 0.05fF
C37 GND a_16444_n18992# 0.02fF
C38 w_15825_n19127# n2 0.03fF
C39 a_16221_n19167# w_16164_n19124# 0.09fF
C40 CompB0 y3 0.11fF
C41 CompB2not y3 0.11fF
C42 y0 y3 0.20fF
C43 a_15955_n19164# VDD 0.12fF
C44 a_16444_n18992# n1 0.08fF
C45 w_16219_n19300# n1 0.08fF
C46 CompB3not a_15514_n19318# 0.17fF
C47 w_16431_n18998# n0 0.08fF
C48 CompB1 w_15942_n19124# 0.13fF
C49 CompA0 CompB0 0.79fF
C50 GND AGB 0.17fF
C51 GND a_15999_n19167# 0.04fF
C52 CompB3 a_15475_n19164# 0.10fF
C53 GND CompB3not 0.12fF
C54 y1 w_16019_n19310# 0.03fF
C55 n2 CompB1not 0.77fF
C56 CompB0 a_16203_n19164# 0.10fF
C57 n2 VDD 0.39fF
C58 CompB3 a_15449_n19164# 0.20fF
C59 CompA1 w_15942_n19124# 0.14fF
C60 w_16082_n19127# a_15981_n19164# 0.06fF
C61 a_16232_n19294# VDD 0.21fF
C62 CompB3 w_15436_n19124# 0.13fF
C63 w_15942_n19124# a_15981_n19164# 0.02fF
C64 w_16480_n19371# y2 0.06fF
C65 a_16444_n18992# VDD 0.17fF
C66 w_16219_n19300# VDD 0.08fF
C67 a_16177_n19164# w_16164_n19124# 0.09fF
C68 a_15514_n19318# y3 0.05fF
C69 a_16221_n19167# CompB0 0.28fF
C70 w_16019_n19310# VDD 0.03fF
C71 GND y3 0.22fF
C72 GND a_15742_n19167# 0.04fF
C73 y0 w_16480_n19371# 0.06fF
C74 AGB VDD 0.16fF
C75 a_15999_n19167# VDD 0.06fF
C76 GND ALB 0.13fF
C77 GND a_15475_n19164# 0.01fF
C78 CompB3not VDD 0.13fF
C79 a_16232_n19294# n2 0.16fF
C80 CompA1 a_15971_n19304# 0.12fF
C81 y0 w_16292_n19300# 0.03fF
C82 n3 a_15971_n19304# 0.04fF
C83 y1 y3 0.20fF
C84 CompB3 CompA3 0.76fF
C85 GND CompA0 0.17fF
C86 n2 a_16444_n18992# 0.16fF
C87 GND a_15449_n19164# 0.08fF
C88 n3 CompA2 0.20fF
C89 CompA0 n1 1.99fF
C90 a_15514_n19318# w_15501_n19324# 0.02fF
C91 n2 w_16219_n19300# 0.08fF
C92 GND n0 0.12fF
C93 GND a_16203_n19164# 0.01fF
C94 n1 n0 1.30fF
C95 w_15544_n19324# y3 0.03fF
C96 CompB1 CompA1 0.87fF
C97 AEB GND 0.17fF
C98 CompB1 n3 0.28fF
C99 CompB3 a_15493_n19167# 0.28fF
C100 a_15742_n19167# w_15685_n19124# 0.09fF
C101 a_16232_n19294# w_16219_n19300# 0.08fF
C102 CompB1 a_15981_n19164# 0.10fF
C103 y3 CompB2 0.07fF
C104 w_16480_n19371# a_16493_n19415# 0.09fF
C105 a_15742_n19167# CompB2 0.28fF
C106 CompB1not y3 0.12fF
C107 a_16177_n19164# CompB0 0.20fF
C108 VDD y3 0.06fF
C109 a_15742_n19167# VDD 0.06fF
C110 CompA1 n3 0.19fF
C111 a_15514_n19318# CompA3 0.04fF
C112 GND a_15698_n19164# 0.08fF
C113 GND a_16221_n19167# 0.04fF
C114 CompB1 y2 0.09fF
C115 CompA1 a_15981_n19164# 0.01fF
C116 GND a_15724_n19164# 0.01fF
C117 CompB2not CompA2 0.93fF
C118 GND CompA3 0.08fF
C119 CompA0 VDD 0.34fF
C120 a_15449_n19164# VDD 0.12fF
C121 CompB0not n3 0.08fF
C122 VDD w_15576_n19127# 0.05fF
C123 VDD n0 0.17fF
C124 CompB2not w_15617_n19485# 0.03fF
C125 y1 w_16480_n19371# 0.06fF
C126 w_16082_n19127# n1 0.03fF
C127 VDD w_15436_n19124# 0.12fF
C128 w_15501_n19324# VDD 0.06fF
C129 AEB VDD 0.17fF
C130 CompB0 w_16164_n19124# 0.13fF
C131 GND a_15493_n19167# 0.04fF
C132 w_16730_n19153# VDD 0.03fF
C133 a_15724_n19164# w_15825_n19127# 0.06fF
C134 n3 w_16431_n18998# 0.08fF
C135 a_15698_n19164# w_15685_n19124# 0.09fF
C136 a_15724_n19164# w_15685_n19124# 0.02fF
C137 CompB0not y2 0.10fF
C138 CompB0 n3 0.11fF
C139 CompA0 n2 0.18fF
C140 CompB2not n3 0.46fF
C141 a_15971_n19304# w_15958_n19310# 0.05fF
C142 a_15698_n19164# CompB2 0.20fF
C143 n2 n0 0.08fF
C144 a_15698_n19164# VDD 0.12fF
C145 a_16221_n19167# VDD 0.06fF
C146 a_15724_n19164# CompB2 0.10fF
C147 CompB0not CompB0 0.02fF
C148 a_16232_n19294# CompA0 0.08fF
C149 GND a_16177_n19164# 0.08fF
C150 w_16480_n19371# VDD 0.06fF
C151 CompA3 VDD 0.23fF
C152 GND a_15971_n19304# 0.02fF
C153 w_16292_n19300# VDD 0.03fF
C154 w_16082_n19127# VDD 0.05fF
C155 CompB0 y2 0.11fF
C156 CompA0 w_16219_n19300# 0.08fF
C157 GND CompA2 0.18fF
C158 y0 y2 0.20fF
C159 y1 a_15971_n19304# 0.05fF
C160 AGB ALB 0.19fF
C161 a_16444_n18992# n0 0.12fF
C162 w_15942_n19124# VDD 0.12fF
C163 a_15493_n19167# VDD 0.06fF
C164 AEB a_16444_n18992# 0.05fF
C165 a_15955_n19164# w_15942_n19124# 0.09fF
C166 CompB1 GND 0.24fF
C167 a_15724_n19164# n2 0.02fF
C168 a_15716_n19313# CompA2 0.12fF
C169 CompB3 w_15561_n19485# 0.06fF
C170 CompA1 w_15958_n19310# 0.08fF
C171 n3 w_15958_n19310# 0.08fF
C172 w_15703_n19319# CompA2 0.08fF
C173 AEB AGB 1.80fF
C174 CompB3not w_15501_n19324# 0.08fF
C175 w_15685_n19124# CompA2 0.14fF
C176 AGB w_16730_n19153# 0.06fF
C177 GND CompA1 0.46fF
C178 GND n3 0.17fF
C179 a_16177_n19164# VDD 0.12fF
C180 CompB1not a_15971_n19304# 0.08fF
C181 a_16232_n19294# w_16292_n19300# 0.08fF
C182 a_15971_n19304# VDD 0.17fF
C183 n3 n1 0.26fF
C184 GND a_15981_n19164# 0.01fF
C185 a_16493_n19415# y2 0.08fF
C186 CompA2 CompB2 0.97fF
C187 a_15981_n19164# n1 0.02fF
C188 GND CompB0not 0.30fF
C189 VDD CompA2 0.32fF
C190 CompB0not n1 0.08fF
C191 a_15716_n19313# n3 0.04fF
C192 w_15756_n19319# y2 0.03fF
C193 n3 w_15703_n19319# 0.08fF
C194 w_15617_n19485# CompB2 0.06fF
C195 CompB0not y1 0.10fF
C196 AGB w_16480_n19371# 0.03fF
C197 CompB1 CompB1not 0.16fF
C198 VDD w_16492_n18998# 0.03fF
C199 CompB1 VDD 0.11fF
C200 y0 a_16493_n19415# 0.38fF
C201 w_15617_n19485# VDD 0.05fF
C202 GND y2 0.25fF
C203 CompB1 w_15814_n19485# 0.06fF
C204 w_16304_n19127# VDD 0.05fF
C205 CompB3not CompA3 0.26fF
C206 a_15449_n19164# a_15475_n19164# 0.12fF
C207 w_16164_n19124# VDD 0.12fF
C208 CompB1 a_15955_n19164# 0.20fF
C209 a_15475_n19164# w_15576_n19127# 0.06fF
C210 n2 a_15971_n19304# 0.16fF
C211 w_16431_n18998# n1 0.08fF
C212 y1 y2 6.45fF
C213 w_15942_n19124# a_15999_n19167# 0.09fF
C214 a_15475_n19164# w_15436_n19124# 0.02fF
C215 GND CompB0 0.33fF
C216 GND CompB2not 0.16fF
C217 GND y0 0.06fF
C218 a_15716_n19313# y2 0.05fF
C219 CompA1 CompB1not 0.80fF
C220 n3 CompB2 0.15fF
C221 CompB0 n1 0.11fF
C222 CompA1 VDD 0.26fF
C223 n3 CompB1not 0.08fF
C224 w_16730_n19153# ALB 0.03fF
C225 CompA0 a_16203_n19164# 0.01fF
C226 n3 VDD 0.45fF
C227 a_15449_n19164# w_15436_n19124# 0.09fF
C228 y1 CompB0 0.11fF
C229 a_16203_n19164# n0 0.02fF
C230 GND CompB3 0.13fF
C231 y0 y1 2.34fF
C232 a_15955_n19164# CompA1 0.08fF
C233 CompB0not w_16077_n19485# 0.03fF
C234 CompB1 n2 0.20fF
C235 CompB2not a_15716_n19313# 0.16fF
C236 CompB0not VDD 0.15fF
C237 CompB2not w_15703_n19319# 0.08fF
C238 a_15955_n19164# a_15981_n19164# 0.12fF
C239 a_15971_n19304# w_16019_n19310# 0.08fF
C240 a_15742_n19167# a_15724_n19164# 0.09fF
C241 w_16480_n19371# y3 0.06fF
C242 AEB w_16730_n19153# 0.06fF
C243 CompB1not y2 0.10fF
C244 VDD y2 0.06fF
C245 CompA3 a_15475_n19164# 0.01fF
C246 CompA1 n2 1.00fF
C247 n3 n2 10.84fF
C248 a_16444_n18992# w_16492_n18998# 0.08fF
C249 VDD w_16431_n18998# 0.08fF
C250 a_16221_n19167# CompA0 0.10fF
C251 w_15561_n19485# VDD 0.05fF
C252 CompB0 w_16077_n19485# 0.06fF
C253 CompB2not CompB2 0.02fF
C254 GND a_16493_n19415# 0.25fF
C255 a_15449_n19164# CompA3 0.08fF
C256 a_16221_n19167# a_16203_n19164# 0.09fF
C257 CompB0 VDD 0.20fF
C258 CompB2not VDD 0.14fF
C259 y0 VDD 0.06fF
C260 CompB0not n2 0.08fF
C261 a_16232_n19294# n3 0.04fF
C262 a_15493_n19167# a_15475_n19164# 0.09fF
C263 GND a_15514_n19318# 0.02fF
C264 CompB1 a_15999_n19167# 0.28fF
C265 y1 a_16493_n19415# 0.08fF
C266 CompA3 w_15436_n19124# 0.14fF
C267 CompA3 w_15501_n19324# 0.08fF
C268 n3 a_16444_n18992# 0.04fF
C269 CompB0not a_16232_n19294# 0.12fF
C270 n3 w_16219_n19300# 0.08fF
C271 GND n1 0.18fF
C272 n2 w_16431_n18998# 0.08fF
C273 a_15716_n19313# w_15756_n19319# 0.08fF
C274 GND y1 0.26fF
C275 a_15493_n19167# w_15436_n19124# 0.09fF
C276 CompA1 a_15999_n19167# 0.10fF
C277 CompB0not w_16219_n19300# 0.08fF
C278 CompB0 n2 0.11fF
C279 GND a_15716_n19313# 0.02fF
C280 a_15698_n19164# a_15724_n19164# 0.12fF
C281 a_15514_n19318# w_15544_n19324# 0.08fF
C282 a_15999_n19167# a_15981_n19164# 0.09fF
C283 a_15742_n19167# CompA2 0.10fF
C284 a_16444_n18992# w_16431_n18998# 0.05fF
C285 a_16177_n19164# CompA0 0.08fF
C286 VDD a_16493_n19415# 0.04fF
C287 a_16232_n19294# y0 0.05fF
C288 CompB1not w_15958_n19310# 0.08fF
C289 w_15958_n19310# VDD 0.08fF
C290 a_16177_n19164# a_16203_n19164# 0.12fF
C291 a_15716_n19313# w_15703_n19319# 0.05fF
C292 CompB1 y3 0.07fF
C293 a_15514_n19318# VDD 0.09fF
C294 w_15756_n19319# VDD 0.03fF
C295 GND CompB2 0.25fF
C296 GND CompB1not 0.18fF
C297 CompA3 a_15493_n19167# 0.10fF
C298 a_16493_n19415# Gnd 0.54fF
C299 y2 Gnd 0.11fF
C300 y1 Gnd 0.14fF
C301 a_15716_n19313# Gnd 0.43fF
C302 CompB2not Gnd 0.06fF
C303 a_15514_n19318# Gnd 0.37fF
C304 CompB3not Gnd 0.25fF
C305 y0 Gnd 2.13fF
C306 a_15971_n19304# Gnd 0.52fF
C307 CompB1not Gnd 0.06fF
C308 a_16232_n19294# Gnd 0.08fF
C309 CompB0not Gnd 0.06fF
C310 ALB Gnd 0.14fF
C311 AGB Gnd 1.78fF
C312 a_16203_n19164# Gnd 1.03fF
C313 a_16221_n19167# Gnd 0.42fF
C314 a_16177_n19164# Gnd 0.50fF
C315 CompB0 Gnd 0.18fF
C316 CompA0 Gnd 4.40fF
C317 a_15981_n19164# Gnd 1.03fF
C318 a_15999_n19167# Gnd 0.42fF
C319 CompB1 Gnd 0.18fF
C320 CompA1 Gnd 0.26fF
C321 a_15724_n19164# Gnd 0.08fF
C322 a_15742_n19167# Gnd 0.21fF
C323 a_15698_n19164# Gnd 0.39fF
C324 CompB2 Gnd 0.32fF
C325 CompA2 Gnd 0.26fF
C326 a_15475_n19164# Gnd 1.03fF
C327 a_15493_n19167# Gnd 0.42fF
C328 a_15449_n19164# Gnd 0.09fF
C329 CompA3 Gnd 0.25fF
C330 GND Gnd 0.09fF
C331 AEB Gnd 1.62fF
C332 VDD Gnd 25.09fF
C333 a_16444_n18992# Gnd 0.03fF
C334 n0 Gnd 0.06fF
C335 n1 Gnd 0.06fF
C336 n2 Gnd 0.06fF
C337 n3 Gnd 0.06fF
C338 w_16077_n19485# Gnd 0.40fF
C339 w_15814_n19485# Gnd 0.40fF
C340 w_15617_n19485# Gnd 0.40fF
C341 w_15561_n19485# Gnd 0.40fF
C342 w_16480_n19371# Gnd 1.36fF
C343 w_16292_n19300# Gnd 0.43fF
C344 w_16219_n19300# Gnd 0.65fF
C345 w_16019_n19310# Gnd 0.43fF
C346 w_15958_n19310# Gnd 0.99fF
C347 w_15756_n19319# Gnd 0.43fF
C348 w_15703_n19319# Gnd 0.83fF
C349 w_15544_n19324# Gnd 0.43fF
C350 w_15501_n19324# Gnd 0.67fF
C351 w_16730_n19153# Gnd 0.45fF
C352 w_16304_n19127# Gnd 0.40fF
C353 w_16164_n19124# Gnd 1.63fF
C354 w_16082_n19127# Gnd 0.40fF
C355 w_15942_n19124# Gnd 1.63fF
C356 w_15825_n19127# Gnd 0.40fF
C357 w_15685_n19124# Gnd 1.63fF
C358 w_15576_n19127# Gnd 0.40fF
C359 w_15436_n19124# Gnd 1.63fF
C360 w_16492_n18998# Gnd 0.43fF
C361 w_16431_n18998# Gnd 0.43fF
.tran 0.05n 100n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(CompA0) v(CompA1)+3 v(CompA2)+6 v(CompA3)+9  v(CompB0)+12 v(CompB1)+15 v(CompB2)+18 v(CompB3)+21 
plot v(ALB) v(AEB)+3 v(AGB)+6

.endc
.end