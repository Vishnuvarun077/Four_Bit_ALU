magic
tech scmos
timestamp 1701461277
<< nwell >>
rect 16431 -18998 16486 -18980
rect 16492 -18998 16516 -18980
rect 15436 -19124 15526 -19106
rect 15576 -19127 15601 -19111
rect 15685 -19124 15775 -19106
rect 15825 -19127 15850 -19111
rect 15942 -19124 16032 -19106
rect 16082 -19127 16107 -19111
rect 16164 -19124 16254 -19106
rect 16304 -19127 16329 -19111
rect 16730 -19153 16764 -19135
rect 15501 -19324 15538 -19306
rect 15544 -19324 15568 -19306
rect 15703 -19319 15749 -19301
rect 15756 -19319 15780 -19301
rect 15958 -19310 16013 -19292
rect 16019 -19310 16043 -19292
rect 16219 -19300 16284 -19282
rect 16292 -19300 16316 -19282
rect 16480 -19371 16557 -19353
rect 15561 -19485 15586 -19469
rect 15617 -19485 15642 -19469
rect 15814 -19485 15839 -19469
rect 16077 -19485 16102 -19469
<< ntransistor >>
rect 16442 -19033 16444 -19029
rect 16452 -19033 16454 -19029
rect 16462 -19033 16464 -19029
rect 16472 -19033 16474 -19029
rect 16503 -19033 16505 -19029
rect 15587 -19141 15589 -19137
rect 15447 -19164 15449 -19160
rect 15463 -19164 15465 -19160
rect 15473 -19164 15475 -19160
rect 15483 -19164 15485 -19160
rect 15493 -19164 15495 -19160
rect 15836 -19141 15838 -19137
rect 15513 -19164 15515 -19160
rect 15696 -19164 15698 -19160
rect 15712 -19164 15714 -19160
rect 15722 -19164 15724 -19160
rect 15732 -19164 15734 -19160
rect 15742 -19164 15744 -19160
rect 16093 -19141 16095 -19137
rect 15762 -19164 15764 -19160
rect 15953 -19164 15955 -19160
rect 15969 -19164 15971 -19160
rect 15979 -19164 15981 -19160
rect 15989 -19164 15991 -19160
rect 15999 -19164 16001 -19160
rect 16315 -19141 16317 -19137
rect 16019 -19164 16021 -19160
rect 16175 -19164 16177 -19160
rect 16191 -19164 16193 -19160
rect 16201 -19164 16203 -19160
rect 16211 -19164 16213 -19160
rect 16221 -19164 16223 -19160
rect 16241 -19164 16243 -19160
rect 16741 -19183 16743 -19179
rect 16751 -19183 16753 -19179
rect 15512 -19348 15514 -19344
rect 15522 -19348 15524 -19344
rect 15555 -19348 15557 -19344
rect 15714 -19346 15716 -19342
rect 15724 -19346 15726 -19342
rect 15734 -19346 15736 -19342
rect 15767 -19346 15769 -19342
rect 15969 -19345 15971 -19341
rect 15979 -19345 15981 -19341
rect 15989 -19345 15991 -19341
rect 15999 -19345 16001 -19341
rect 16030 -19345 16032 -19341
rect 16230 -19342 16232 -19338
rect 16240 -19342 16242 -19338
rect 16250 -19342 16252 -19338
rect 16260 -19342 16262 -19338
rect 16270 -19342 16272 -19338
rect 16303 -19342 16305 -19338
rect 16491 -19415 16493 -19411
rect 16501 -19415 16503 -19411
rect 16510 -19415 16512 -19411
rect 16520 -19415 16522 -19411
rect 16539 -19415 16541 -19411
rect 15572 -19499 15574 -19495
rect 15628 -19499 15630 -19495
rect 15825 -19499 15827 -19495
rect 16088 -19499 16090 -19495
<< ptransistor >>
rect 16442 -18992 16444 -18986
rect 16452 -18992 16454 -18986
rect 16462 -18992 16464 -18986
rect 16472 -18992 16474 -18986
rect 16503 -18992 16505 -18986
rect 15447 -19118 15449 -19112
rect 15463 -19118 15465 -19112
rect 15473 -19118 15475 -19112
rect 15483 -19118 15485 -19112
rect 15493 -19118 15495 -19112
rect 15513 -19118 15515 -19112
rect 15587 -19121 15589 -19117
rect 15696 -19118 15698 -19112
rect 15712 -19118 15714 -19112
rect 15722 -19118 15724 -19112
rect 15732 -19118 15734 -19112
rect 15742 -19118 15744 -19112
rect 15762 -19118 15764 -19112
rect 15836 -19121 15838 -19117
rect 15953 -19118 15955 -19112
rect 15969 -19118 15971 -19112
rect 15979 -19118 15981 -19112
rect 15989 -19118 15991 -19112
rect 15999 -19118 16001 -19112
rect 16019 -19118 16021 -19112
rect 16093 -19121 16095 -19117
rect 16175 -19118 16177 -19112
rect 16191 -19118 16193 -19112
rect 16201 -19118 16203 -19112
rect 16211 -19118 16213 -19112
rect 16221 -19118 16223 -19112
rect 16241 -19118 16243 -19112
rect 16315 -19121 16317 -19117
rect 16741 -19147 16743 -19141
rect 16751 -19147 16753 -19141
rect 16230 -19294 16232 -19288
rect 16240 -19294 16242 -19288
rect 16250 -19294 16252 -19288
rect 16260 -19294 16262 -19288
rect 16270 -19294 16272 -19288
rect 16303 -19294 16305 -19288
rect 15969 -19304 15971 -19298
rect 15979 -19304 15981 -19298
rect 15989 -19304 15991 -19298
rect 15999 -19304 16001 -19298
rect 16030 -19304 16032 -19298
rect 15512 -19318 15514 -19312
rect 15522 -19318 15524 -19312
rect 15555 -19318 15557 -19312
rect 15714 -19313 15716 -19307
rect 15724 -19313 15726 -19307
rect 15734 -19313 15736 -19307
rect 15767 -19313 15769 -19307
rect 16491 -19365 16493 -19359
rect 16501 -19365 16503 -19359
rect 16510 -19365 16512 -19359
rect 16520 -19365 16522 -19359
rect 16539 -19365 16541 -19359
rect 15572 -19479 15574 -19475
rect 15628 -19479 15630 -19475
rect 15825 -19479 15827 -19475
rect 16088 -19479 16090 -19475
<< ndiffusion >>
rect 16441 -19033 16442 -19029
rect 16444 -19033 16452 -19029
rect 16454 -19033 16462 -19029
rect 16464 -19033 16472 -19029
rect 16474 -19033 16476 -19029
rect 16502 -19033 16503 -19029
rect 16505 -19033 16506 -19029
rect 15586 -19141 15587 -19137
rect 15589 -19141 15590 -19137
rect 15446 -19164 15447 -19160
rect 15449 -19164 15450 -19160
rect 15462 -19164 15463 -19160
rect 15465 -19164 15473 -19160
rect 15475 -19164 15477 -19160
rect 15481 -19164 15483 -19160
rect 15485 -19164 15493 -19160
rect 15495 -19164 15496 -19160
rect 15835 -19141 15836 -19137
rect 15838 -19141 15839 -19137
rect 15512 -19164 15513 -19160
rect 15515 -19164 15516 -19160
rect 15695 -19164 15696 -19160
rect 15698 -19164 15699 -19160
rect 15711 -19164 15712 -19160
rect 15714 -19164 15722 -19160
rect 15724 -19164 15726 -19160
rect 15730 -19164 15732 -19160
rect 15734 -19164 15742 -19160
rect 15744 -19164 15745 -19160
rect 16092 -19141 16093 -19137
rect 16095 -19141 16096 -19137
rect 15761 -19164 15762 -19160
rect 15764 -19164 15765 -19160
rect 15952 -19164 15953 -19160
rect 15955 -19164 15956 -19160
rect 15968 -19164 15969 -19160
rect 15971 -19164 15979 -19160
rect 15981 -19164 15983 -19160
rect 15987 -19164 15989 -19160
rect 15991 -19164 15999 -19160
rect 16001 -19164 16002 -19160
rect 16314 -19141 16315 -19137
rect 16317 -19141 16318 -19137
rect 16018 -19164 16019 -19160
rect 16021 -19164 16022 -19160
rect 16174 -19164 16175 -19160
rect 16177 -19164 16178 -19160
rect 16190 -19164 16191 -19160
rect 16193 -19164 16201 -19160
rect 16203 -19164 16205 -19160
rect 16209 -19164 16211 -19160
rect 16213 -19164 16221 -19160
rect 16223 -19164 16224 -19160
rect 16240 -19164 16241 -19160
rect 16243 -19164 16244 -19160
rect 16740 -19183 16741 -19179
rect 16743 -19183 16745 -19179
rect 16749 -19183 16751 -19179
rect 16753 -19183 16754 -19179
rect 15511 -19348 15512 -19344
rect 15514 -19348 15522 -19344
rect 15524 -19348 15526 -19344
rect 15554 -19348 15555 -19344
rect 15557 -19348 15558 -19344
rect 15713 -19346 15714 -19342
rect 15716 -19346 15724 -19342
rect 15726 -19346 15734 -19342
rect 15736 -19346 15738 -19342
rect 15766 -19346 15767 -19342
rect 15769 -19346 15770 -19342
rect 15968 -19345 15969 -19341
rect 15971 -19345 15979 -19341
rect 15981 -19345 15989 -19341
rect 15991 -19345 15999 -19341
rect 16001 -19345 16003 -19341
rect 16029 -19345 16030 -19341
rect 16032 -19345 16033 -19341
rect 16229 -19342 16230 -19338
rect 16232 -19342 16240 -19338
rect 16242 -19342 16250 -19338
rect 16252 -19342 16260 -19338
rect 16262 -19342 16270 -19338
rect 16272 -19342 16274 -19338
rect 16302 -19342 16303 -19338
rect 16305 -19342 16306 -19338
rect 16490 -19415 16491 -19411
rect 16493 -19415 16495 -19411
rect 16499 -19415 16501 -19411
rect 16503 -19415 16504 -19411
rect 16508 -19415 16510 -19411
rect 16512 -19415 16514 -19411
rect 16518 -19415 16520 -19411
rect 16522 -19415 16524 -19411
rect 16538 -19415 16539 -19411
rect 16541 -19415 16542 -19411
rect 15571 -19499 15572 -19495
rect 15574 -19499 15575 -19495
rect 15627 -19499 15628 -19495
rect 15630 -19499 15631 -19495
rect 15824 -19499 15825 -19495
rect 15827 -19499 15828 -19495
rect 16087 -19499 16088 -19495
rect 16090 -19499 16091 -19495
<< pdiffusion >>
rect 16441 -18992 16442 -18986
rect 16444 -18992 16446 -18986
rect 16450 -18992 16452 -18986
rect 16454 -18992 16456 -18986
rect 16460 -18992 16462 -18986
rect 16464 -18992 16466 -18986
rect 16470 -18992 16472 -18986
rect 16474 -18992 16476 -18986
rect 16502 -18992 16503 -18986
rect 16505 -18992 16506 -18986
rect 15446 -19118 15447 -19112
rect 15449 -19118 15450 -19112
rect 15462 -19118 15463 -19112
rect 15465 -19118 15473 -19112
rect 15475 -19118 15477 -19112
rect 15481 -19118 15483 -19112
rect 15485 -19118 15493 -19112
rect 15495 -19118 15496 -19112
rect 15512 -19118 15513 -19112
rect 15515 -19118 15516 -19112
rect 15586 -19121 15587 -19117
rect 15589 -19121 15590 -19117
rect 15695 -19118 15696 -19112
rect 15698 -19118 15699 -19112
rect 15711 -19118 15712 -19112
rect 15714 -19118 15722 -19112
rect 15724 -19118 15726 -19112
rect 15730 -19118 15732 -19112
rect 15734 -19118 15742 -19112
rect 15744 -19118 15745 -19112
rect 15761 -19118 15762 -19112
rect 15764 -19118 15765 -19112
rect 15835 -19121 15836 -19117
rect 15838 -19121 15839 -19117
rect 15952 -19118 15953 -19112
rect 15955 -19118 15956 -19112
rect 15968 -19118 15969 -19112
rect 15971 -19118 15979 -19112
rect 15981 -19118 15983 -19112
rect 15987 -19118 15989 -19112
rect 15991 -19118 15999 -19112
rect 16001 -19118 16002 -19112
rect 16018 -19118 16019 -19112
rect 16021 -19118 16022 -19112
rect 16092 -19121 16093 -19117
rect 16095 -19121 16096 -19117
rect 16174 -19118 16175 -19112
rect 16177 -19118 16178 -19112
rect 16190 -19118 16191 -19112
rect 16193 -19118 16201 -19112
rect 16203 -19118 16205 -19112
rect 16209 -19118 16211 -19112
rect 16213 -19118 16221 -19112
rect 16223 -19118 16224 -19112
rect 16240 -19118 16241 -19112
rect 16243 -19118 16244 -19112
rect 16314 -19121 16315 -19117
rect 16317 -19121 16318 -19117
rect 16740 -19147 16741 -19141
rect 16743 -19147 16751 -19141
rect 16753 -19147 16754 -19141
rect 16229 -19294 16230 -19288
rect 16232 -19294 16234 -19288
rect 16238 -19294 16240 -19288
rect 16242 -19294 16244 -19288
rect 16248 -19294 16250 -19288
rect 16252 -19294 16254 -19288
rect 16258 -19294 16260 -19288
rect 16262 -19294 16264 -19288
rect 16268 -19294 16270 -19288
rect 16272 -19294 16274 -19288
rect 16302 -19294 16303 -19288
rect 16305 -19294 16306 -19288
rect 15968 -19304 15969 -19298
rect 15971 -19304 15973 -19298
rect 15977 -19304 15979 -19298
rect 15981 -19304 15983 -19298
rect 15987 -19304 15989 -19298
rect 15991 -19304 15993 -19298
rect 15997 -19304 15999 -19298
rect 16001 -19304 16003 -19298
rect 16029 -19304 16030 -19298
rect 16032 -19304 16033 -19298
rect 15511 -19318 15512 -19312
rect 15514 -19318 15516 -19312
rect 15520 -19318 15522 -19312
rect 15524 -19318 15526 -19312
rect 15554 -19318 15555 -19312
rect 15557 -19318 15558 -19312
rect 15713 -19313 15714 -19307
rect 15716 -19313 15718 -19307
rect 15722 -19313 15724 -19307
rect 15726 -19313 15728 -19307
rect 15732 -19313 15734 -19307
rect 15736 -19313 15738 -19307
rect 15766 -19313 15767 -19307
rect 15769 -19313 15770 -19307
rect 16490 -19365 16491 -19359
rect 16493 -19365 16501 -19359
rect 16503 -19365 16510 -19359
rect 16512 -19365 16520 -19359
rect 16522 -19365 16524 -19359
rect 16538 -19365 16539 -19359
rect 16541 -19365 16542 -19359
rect 15571 -19479 15572 -19475
rect 15574 -19479 15575 -19475
rect 15627 -19479 15628 -19475
rect 15630 -19479 15631 -19475
rect 15824 -19479 15825 -19475
rect 15827 -19479 15828 -19475
rect 16087 -19479 16088 -19475
rect 16090 -19479 16091 -19475
<< ndcontact >>
rect 16437 -19033 16441 -19029
rect 16476 -19033 16480 -19029
rect 16498 -19033 16502 -19029
rect 16506 -19033 16510 -19029
rect 15582 -19141 15586 -19137
rect 15590 -19141 15594 -19137
rect 15442 -19164 15446 -19160
rect 15450 -19164 15454 -19160
rect 15458 -19164 15462 -19160
rect 15477 -19164 15481 -19160
rect 15496 -19164 15500 -19160
rect 15831 -19141 15835 -19137
rect 15839 -19141 15843 -19137
rect 15508 -19164 15512 -19160
rect 15516 -19164 15520 -19160
rect 15691 -19164 15695 -19160
rect 15699 -19164 15703 -19160
rect 15707 -19164 15711 -19160
rect 15726 -19164 15730 -19160
rect 15745 -19164 15749 -19160
rect 16088 -19141 16092 -19137
rect 16096 -19141 16100 -19137
rect 15757 -19164 15761 -19160
rect 15765 -19164 15769 -19160
rect 15948 -19164 15952 -19160
rect 15956 -19164 15960 -19160
rect 15964 -19164 15968 -19160
rect 15983 -19164 15987 -19160
rect 16002 -19164 16006 -19160
rect 16310 -19141 16314 -19137
rect 16318 -19141 16322 -19137
rect 16014 -19164 16018 -19160
rect 16022 -19164 16026 -19160
rect 16170 -19164 16174 -19160
rect 16178 -19164 16182 -19160
rect 16186 -19164 16190 -19160
rect 16205 -19164 16209 -19160
rect 16224 -19164 16228 -19160
rect 16236 -19164 16240 -19160
rect 16244 -19164 16248 -19160
rect 16736 -19183 16740 -19179
rect 16745 -19183 16749 -19179
rect 16754 -19183 16758 -19179
rect 15507 -19348 15511 -19344
rect 15526 -19348 15530 -19344
rect 15550 -19348 15554 -19344
rect 15558 -19348 15562 -19344
rect 15709 -19346 15713 -19342
rect 15738 -19346 15742 -19342
rect 15762 -19346 15766 -19342
rect 15770 -19346 15774 -19342
rect 15964 -19345 15968 -19341
rect 16003 -19345 16007 -19341
rect 16025 -19345 16029 -19341
rect 16033 -19345 16037 -19341
rect 16225 -19342 16229 -19338
rect 16274 -19342 16278 -19338
rect 16298 -19342 16302 -19338
rect 16306 -19342 16310 -19338
rect 16486 -19415 16490 -19411
rect 16495 -19415 16499 -19411
rect 16504 -19415 16508 -19411
rect 16514 -19415 16518 -19411
rect 16524 -19415 16528 -19411
rect 16534 -19415 16538 -19411
rect 16542 -19415 16546 -19411
rect 15567 -19499 15571 -19495
rect 15575 -19499 15579 -19495
rect 15623 -19499 15627 -19495
rect 15631 -19499 15635 -19495
rect 15820 -19499 15824 -19495
rect 15828 -19499 15832 -19495
rect 16083 -19499 16087 -19495
rect 16091 -19499 16095 -19495
<< pdcontact >>
rect 16437 -18992 16441 -18986
rect 16446 -18992 16450 -18986
rect 16456 -18992 16460 -18986
rect 16466 -18992 16470 -18986
rect 16476 -18992 16480 -18986
rect 16498 -18992 16502 -18986
rect 16506 -18992 16510 -18986
rect 15442 -19118 15446 -19112
rect 15450 -19118 15454 -19112
rect 15458 -19118 15462 -19112
rect 15477 -19118 15481 -19112
rect 15496 -19118 15500 -19112
rect 15508 -19118 15512 -19112
rect 15516 -19118 15520 -19112
rect 15582 -19121 15586 -19117
rect 15590 -19121 15594 -19117
rect 15691 -19118 15695 -19112
rect 15699 -19118 15703 -19112
rect 15707 -19118 15711 -19112
rect 15726 -19118 15730 -19112
rect 15745 -19118 15749 -19112
rect 15757 -19118 15761 -19112
rect 15765 -19118 15769 -19112
rect 15831 -19121 15835 -19117
rect 15839 -19121 15843 -19117
rect 15948 -19118 15952 -19112
rect 15956 -19118 15960 -19112
rect 15964 -19118 15968 -19112
rect 15983 -19118 15987 -19112
rect 16002 -19118 16006 -19112
rect 16014 -19118 16018 -19112
rect 16022 -19118 16026 -19112
rect 16088 -19121 16092 -19117
rect 16096 -19121 16100 -19117
rect 16170 -19118 16174 -19112
rect 16178 -19118 16182 -19112
rect 16186 -19118 16190 -19112
rect 16205 -19118 16209 -19112
rect 16224 -19118 16228 -19112
rect 16236 -19118 16240 -19112
rect 16244 -19118 16248 -19112
rect 16310 -19121 16314 -19117
rect 16318 -19121 16322 -19117
rect 16736 -19147 16740 -19141
rect 16754 -19147 16758 -19141
rect 16225 -19294 16229 -19288
rect 16234 -19294 16238 -19288
rect 16244 -19294 16248 -19288
rect 16254 -19294 16258 -19288
rect 16264 -19294 16268 -19288
rect 16274 -19294 16278 -19288
rect 16298 -19294 16302 -19288
rect 16306 -19294 16310 -19288
rect 15964 -19304 15968 -19298
rect 15973 -19304 15977 -19298
rect 15983 -19304 15987 -19298
rect 15993 -19304 15997 -19298
rect 16003 -19304 16007 -19298
rect 16025 -19304 16029 -19298
rect 16033 -19304 16037 -19298
rect 15507 -19318 15511 -19312
rect 15516 -19318 15520 -19312
rect 15526 -19318 15530 -19312
rect 15550 -19318 15554 -19312
rect 15558 -19318 15562 -19312
rect 15709 -19313 15713 -19307
rect 15718 -19313 15722 -19307
rect 15728 -19313 15732 -19307
rect 15738 -19313 15742 -19307
rect 15762 -19313 15766 -19307
rect 15770 -19313 15774 -19307
rect 16486 -19365 16490 -19359
rect 16524 -19365 16528 -19359
rect 16534 -19365 16538 -19359
rect 16542 -19365 16546 -19359
rect 15567 -19479 15571 -19475
rect 15575 -19479 15579 -19475
rect 15623 -19479 15627 -19475
rect 15631 -19479 15635 -19475
rect 15820 -19479 15824 -19475
rect 15828 -19479 15832 -19475
rect 16083 -19479 16087 -19475
rect 16091 -19479 16095 -19475
<< polysilicon >>
rect 16442 -18986 16444 -18977
rect 16452 -18986 16454 -18977
rect 16462 -18986 16464 -18977
rect 16472 -18986 16474 -18977
rect 16503 -18986 16505 -18977
rect 16442 -19029 16444 -18992
rect 16452 -19029 16454 -18992
rect 16462 -19029 16464 -18992
rect 16472 -19029 16474 -18992
rect 16503 -19029 16505 -18992
rect 16442 -19036 16444 -19033
rect 16452 -19036 16454 -19033
rect 16462 -19036 16464 -19033
rect 16472 -19036 16474 -19033
rect 16503 -19036 16505 -19033
rect 15447 -19104 15533 -19102
rect 15447 -19112 15449 -19104
rect 15463 -19112 15465 -19109
rect 15473 -19112 15475 -19109
rect 15483 -19112 15485 -19104
rect 15493 -19112 15495 -19109
rect 15513 -19112 15515 -19109
rect 15447 -19160 15449 -19118
rect 15463 -19160 15465 -19118
rect 15473 -19139 15475 -19118
rect 15483 -19121 15485 -19118
rect 15473 -19141 15485 -19139
rect 15473 -19160 15475 -19157
rect 15483 -19160 15485 -19141
rect 15493 -19160 15495 -19118
rect 15513 -19141 15515 -19118
rect 15531 -19146 15533 -19104
rect 15696 -19104 15782 -19102
rect 15696 -19112 15698 -19104
rect 15712 -19112 15714 -19109
rect 15722 -19112 15724 -19109
rect 15732 -19112 15734 -19104
rect 15742 -19112 15744 -19109
rect 15762 -19112 15764 -19109
rect 15587 -19117 15589 -19114
rect 15587 -19130 15589 -19121
rect 15583 -19132 15589 -19130
rect 15587 -19137 15589 -19132
rect 15587 -19144 15589 -19141
rect 15504 -19148 15533 -19146
rect 15447 -19167 15449 -19164
rect 15463 -19175 15465 -19164
rect 15473 -19170 15475 -19164
rect 15483 -19167 15485 -19164
rect 15493 -19167 15495 -19164
rect 15504 -19170 15506 -19148
rect 15513 -19160 15515 -19152
rect 15696 -19160 15698 -19118
rect 15712 -19160 15714 -19118
rect 15722 -19139 15724 -19118
rect 15732 -19121 15734 -19118
rect 15722 -19141 15734 -19139
rect 15722 -19160 15724 -19157
rect 15732 -19160 15734 -19141
rect 15742 -19160 15744 -19118
rect 15762 -19141 15764 -19118
rect 15780 -19146 15782 -19104
rect 15953 -19104 16039 -19102
rect 15953 -19112 15955 -19104
rect 15969 -19112 15971 -19109
rect 15979 -19112 15981 -19109
rect 15989 -19112 15991 -19104
rect 15999 -19112 16001 -19109
rect 16019 -19112 16021 -19109
rect 15836 -19117 15838 -19114
rect 15836 -19130 15838 -19121
rect 15832 -19132 15838 -19130
rect 15836 -19137 15838 -19132
rect 15836 -19144 15838 -19141
rect 15753 -19148 15782 -19146
rect 15473 -19172 15506 -19170
rect 15513 -19175 15515 -19164
rect 15696 -19167 15698 -19164
rect 15463 -19177 15515 -19175
rect 15712 -19175 15714 -19164
rect 15722 -19170 15724 -19164
rect 15732 -19167 15734 -19164
rect 15742 -19167 15744 -19164
rect 15753 -19170 15755 -19148
rect 15762 -19160 15764 -19152
rect 15953 -19160 15955 -19118
rect 15969 -19160 15971 -19118
rect 15979 -19139 15981 -19118
rect 15989 -19121 15991 -19118
rect 15979 -19141 15991 -19139
rect 15979 -19160 15981 -19157
rect 15989 -19160 15991 -19141
rect 15999 -19160 16001 -19118
rect 16019 -19141 16021 -19118
rect 16037 -19146 16039 -19104
rect 16175 -19104 16261 -19102
rect 16175 -19112 16177 -19104
rect 16191 -19112 16193 -19109
rect 16201 -19112 16203 -19109
rect 16211 -19112 16213 -19104
rect 16221 -19112 16223 -19109
rect 16241 -19112 16243 -19109
rect 16093 -19117 16095 -19114
rect 16093 -19130 16095 -19121
rect 16089 -19132 16095 -19130
rect 16093 -19137 16095 -19132
rect 16093 -19144 16095 -19141
rect 16010 -19148 16039 -19146
rect 15722 -19172 15755 -19170
rect 15762 -19175 15764 -19164
rect 15953 -19167 15955 -19164
rect 15712 -19177 15764 -19175
rect 15969 -19175 15971 -19164
rect 15979 -19170 15981 -19164
rect 15989 -19167 15991 -19164
rect 15999 -19167 16001 -19164
rect 16010 -19170 16012 -19148
rect 16019 -19160 16021 -19152
rect 16175 -19160 16177 -19118
rect 16191 -19160 16193 -19118
rect 16201 -19139 16203 -19118
rect 16211 -19121 16213 -19118
rect 16201 -19141 16213 -19139
rect 16201 -19160 16203 -19157
rect 16211 -19160 16213 -19141
rect 16221 -19160 16223 -19118
rect 16241 -19141 16243 -19118
rect 16259 -19146 16261 -19104
rect 16315 -19117 16317 -19114
rect 16315 -19130 16317 -19121
rect 16311 -19132 16317 -19130
rect 16315 -19137 16317 -19132
rect 16741 -19141 16743 -19138
rect 16751 -19141 16753 -19138
rect 16315 -19144 16317 -19141
rect 16232 -19148 16261 -19146
rect 15979 -19172 16012 -19170
rect 16019 -19175 16021 -19164
rect 16175 -19167 16177 -19164
rect 15969 -19177 16021 -19175
rect 16191 -19175 16193 -19164
rect 16201 -19170 16203 -19164
rect 16211 -19167 16213 -19164
rect 16221 -19167 16223 -19164
rect 16232 -19170 16234 -19148
rect 16241 -19160 16243 -19152
rect 16201 -19172 16234 -19170
rect 16241 -19175 16243 -19164
rect 16191 -19177 16243 -19175
rect 16741 -19179 16743 -19147
rect 16751 -19179 16753 -19147
rect 16741 -19186 16743 -19183
rect 16751 -19186 16753 -19183
rect 16230 -19288 16232 -19279
rect 16240 -19288 16242 -19279
rect 16250 -19288 16252 -19279
rect 16260 -19288 16262 -19279
rect 16270 -19288 16272 -19279
rect 16303 -19288 16305 -19279
rect 15969 -19298 15971 -19289
rect 15979 -19298 15981 -19289
rect 15989 -19298 15991 -19289
rect 15999 -19298 16001 -19289
rect 16030 -19298 16032 -19289
rect 15512 -19312 15514 -19303
rect 15522 -19312 15524 -19303
rect 15555 -19312 15557 -19303
rect 15714 -19307 15716 -19298
rect 15724 -19307 15726 -19298
rect 15734 -19307 15736 -19298
rect 15767 -19307 15769 -19298
rect 15512 -19344 15514 -19318
rect 15522 -19344 15524 -19318
rect 15555 -19344 15557 -19318
rect 15714 -19342 15716 -19313
rect 15724 -19342 15726 -19313
rect 15734 -19342 15736 -19313
rect 15767 -19342 15769 -19313
rect 15969 -19341 15971 -19304
rect 15979 -19341 15981 -19304
rect 15989 -19341 15991 -19304
rect 15999 -19341 16001 -19304
rect 16030 -19341 16032 -19304
rect 16230 -19338 16232 -19294
rect 16240 -19338 16242 -19294
rect 16250 -19338 16252 -19294
rect 16260 -19338 16262 -19294
rect 16270 -19338 16272 -19294
rect 16303 -19338 16305 -19294
rect 16230 -19345 16232 -19342
rect 16240 -19345 16242 -19342
rect 16250 -19345 16252 -19342
rect 16260 -19345 16262 -19342
rect 16270 -19345 16272 -19342
rect 16303 -19345 16305 -19342
rect 15512 -19351 15514 -19348
rect 15522 -19351 15524 -19348
rect 15555 -19351 15557 -19348
rect 15714 -19349 15716 -19346
rect 15724 -19349 15726 -19346
rect 15734 -19349 15736 -19346
rect 15767 -19349 15769 -19346
rect 15969 -19348 15971 -19345
rect 15979 -19348 15981 -19345
rect 15989 -19348 15991 -19345
rect 15999 -19348 16001 -19345
rect 16030 -19348 16032 -19345
rect 16491 -19359 16493 -19356
rect 16501 -19359 16503 -19356
rect 16510 -19359 16512 -19356
rect 16520 -19359 16522 -19356
rect 16539 -19359 16541 -19356
rect 16491 -19411 16493 -19365
rect 16501 -19411 16503 -19365
rect 16510 -19388 16512 -19365
rect 16511 -19392 16512 -19388
rect 16510 -19411 16512 -19392
rect 16520 -19411 16522 -19365
rect 16539 -19411 16541 -19365
rect 16491 -19418 16493 -19415
rect 16501 -19418 16503 -19415
rect 16510 -19418 16512 -19415
rect 16520 -19418 16522 -19415
rect 16539 -19418 16541 -19415
rect 15572 -19475 15574 -19472
rect 15628 -19475 15630 -19472
rect 15825 -19475 15827 -19472
rect 16088 -19475 16090 -19472
rect 15572 -19488 15574 -19479
rect 15568 -19490 15574 -19488
rect 15572 -19495 15574 -19490
rect 15628 -19488 15630 -19479
rect 15624 -19490 15630 -19488
rect 15628 -19495 15630 -19490
rect 15825 -19488 15827 -19479
rect 15821 -19490 15827 -19488
rect 15825 -19495 15827 -19490
rect 16088 -19488 16090 -19479
rect 16084 -19490 16090 -19488
rect 16088 -19495 16090 -19490
rect 15572 -19502 15574 -19499
rect 15628 -19502 15630 -19499
rect 15825 -19502 15827 -19499
rect 16088 -19502 16090 -19499
<< polycontact >>
rect 16438 -19004 16442 -19000
rect 16448 -19011 16452 -19007
rect 16458 -19018 16462 -19014
rect 16468 -19025 16472 -19021
rect 16499 -19004 16503 -19000
rect 15443 -19141 15447 -19137
rect 15469 -19141 15473 -19137
rect 15495 -19141 15499 -19137
rect 15515 -19141 15519 -19137
rect 15579 -19133 15583 -19129
rect 15692 -19141 15696 -19137
rect 15515 -19156 15519 -19152
rect 15718 -19141 15722 -19137
rect 15744 -19141 15748 -19137
rect 15764 -19141 15768 -19137
rect 15828 -19133 15832 -19129
rect 15949 -19141 15953 -19137
rect 15764 -19156 15768 -19152
rect 15975 -19141 15979 -19137
rect 16001 -19141 16005 -19137
rect 16021 -19141 16025 -19137
rect 16085 -19133 16089 -19129
rect 16171 -19141 16175 -19137
rect 16021 -19156 16025 -19152
rect 16197 -19141 16201 -19137
rect 16223 -19141 16227 -19137
rect 16243 -19141 16247 -19137
rect 16307 -19133 16311 -19129
rect 16243 -19156 16247 -19152
rect 16737 -19160 16741 -19156
rect 16747 -19167 16751 -19163
rect 15508 -19330 15512 -19326
rect 15518 -19339 15522 -19335
rect 15551 -19330 15555 -19326
rect 15710 -19325 15714 -19321
rect 15720 -19332 15724 -19328
rect 15730 -19339 15734 -19335
rect 15763 -19325 15767 -19321
rect 15965 -19316 15969 -19312
rect 15975 -19323 15979 -19319
rect 15985 -19330 15989 -19326
rect 15995 -19337 15999 -19333
rect 16026 -19316 16030 -19312
rect 16226 -19306 16230 -19302
rect 16236 -19313 16240 -19309
rect 16246 -19320 16250 -19316
rect 16256 -19327 16260 -19323
rect 16266 -19335 16270 -19331
rect 16299 -19306 16303 -19302
rect 16487 -19378 16491 -19374
rect 16497 -19385 16501 -19381
rect 16507 -19392 16511 -19388
rect 16516 -19399 16520 -19395
rect 16535 -19383 16539 -19379
rect 15564 -19491 15568 -19487
rect 15620 -19491 15624 -19487
rect 15817 -19491 15821 -19487
rect 16080 -19491 16084 -19487
<< metal1 >>
rect 16431 -18971 16809 -18967
rect 16437 -18986 16441 -18971
rect 16456 -18986 16460 -18971
rect 16476 -18986 16480 -18971
rect 16498 -18986 16502 -18971
rect 16446 -19000 16450 -18992
rect 16466 -19000 16470 -18992
rect 16506 -19000 16510 -18992
rect 15634 -19004 16438 -19000
rect 16446 -19004 16499 -19000
rect 16506 -19004 16622 -19000
rect 15882 -19011 16448 -19007
rect 16127 -19018 16458 -19014
rect 16375 -19025 16468 -19021
rect 15355 -19084 15423 -19077
rect 15356 -19487 15363 -19084
rect 15436 -19099 16303 -19095
rect 15442 -19112 15446 -19099
rect 15458 -19112 15462 -19099
rect 15496 -19112 15500 -19099
rect 15516 -19112 15520 -19099
rect 15576 -19108 15579 -19099
rect 15576 -19111 15601 -19108
rect 15583 -19117 15586 -19111
rect 15691 -19112 15695 -19099
rect 15707 -19112 15711 -19099
rect 15745 -19112 15749 -19099
rect 15765 -19112 15769 -19099
rect 15825 -19108 15828 -19099
rect 15825 -19111 15850 -19108
rect 15450 -19137 15454 -19118
rect 15477 -19128 15481 -19118
rect 15400 -19141 15443 -19137
rect 15450 -19141 15469 -19137
rect 15400 -19316 15406 -19141
rect 15429 -19149 15436 -19145
rect 15429 -19150 15433 -19149
rect 15450 -19160 15454 -19141
rect 15477 -19160 15481 -19133
rect 15508 -19137 15512 -19118
rect 15832 -19117 15835 -19111
rect 15948 -19112 15952 -19099
rect 15964 -19112 15968 -19099
rect 16002 -19112 16006 -19099
rect 16022 -19112 16026 -19099
rect 16082 -19108 16085 -19099
rect 16082 -19111 16107 -19108
rect 15543 -19133 15579 -19129
rect 15590 -19130 15593 -19121
rect 15590 -19133 15627 -19130
rect 15590 -19137 15593 -19133
rect 15699 -19137 15703 -19118
rect 15726 -19128 15730 -19118
rect 15499 -19141 15512 -19137
rect 15508 -19160 15512 -19141
rect 15519 -19144 15523 -19137
rect 15583 -19145 15586 -19141
rect 15650 -19141 15692 -19137
rect 15699 -19141 15718 -19137
rect 15519 -19156 15523 -19149
rect 15576 -19148 15606 -19145
rect 15442 -19178 15446 -19164
rect 15458 -19178 15462 -19164
rect 15496 -19178 15500 -19164
rect 15516 -19178 15520 -19164
rect 15576 -19178 15579 -19148
rect 15660 -19149 15685 -19145
rect 15699 -19160 15703 -19141
rect 15726 -19160 15730 -19133
rect 15757 -19137 15761 -19118
rect 16089 -19117 16092 -19111
rect 16170 -19112 16174 -19099
rect 16186 -19112 16190 -19099
rect 16224 -19112 16228 -19099
rect 16244 -19112 16248 -19099
rect 16304 -19108 16307 -19099
rect 16304 -19111 16329 -19108
rect 15792 -19133 15828 -19129
rect 15839 -19130 15842 -19121
rect 15839 -19133 15876 -19130
rect 15839 -19137 15842 -19133
rect 15956 -19137 15960 -19118
rect 15983 -19128 15987 -19118
rect 15748 -19141 15761 -19137
rect 15757 -19160 15761 -19141
rect 15768 -19144 15772 -19137
rect 15832 -19145 15835 -19141
rect 15926 -19141 15949 -19137
rect 15956 -19141 15975 -19137
rect 15768 -19156 15772 -19149
rect 15825 -19148 15850 -19145
rect 15691 -19178 15695 -19164
rect 15707 -19178 15711 -19164
rect 15745 -19178 15749 -19164
rect 15765 -19178 15769 -19164
rect 15825 -19178 15828 -19148
rect 15902 -19149 15942 -19145
rect 15956 -19160 15960 -19141
rect 15983 -19160 15987 -19133
rect 16014 -19137 16018 -19118
rect 16311 -19117 16314 -19111
rect 16049 -19133 16085 -19129
rect 16096 -19130 16099 -19121
rect 16096 -19133 16120 -19130
rect 16096 -19137 16099 -19133
rect 16178 -19137 16182 -19118
rect 16205 -19128 16209 -19118
rect 16005 -19141 16018 -19137
rect 16014 -19160 16018 -19141
rect 16025 -19144 16029 -19137
rect 16089 -19145 16092 -19141
rect 16146 -19141 16171 -19137
rect 16178 -19141 16197 -19137
rect 16025 -19156 16029 -19149
rect 16082 -19148 16107 -19145
rect 15948 -19178 15952 -19164
rect 15964 -19178 15968 -19164
rect 16002 -19178 16006 -19164
rect 16022 -19178 16026 -19164
rect 16082 -19178 16085 -19148
rect 16160 -19149 16164 -19145
rect 16178 -19160 16182 -19141
rect 16205 -19160 16209 -19133
rect 16236 -19137 16240 -19118
rect 16271 -19133 16307 -19129
rect 16318 -19130 16321 -19121
rect 16375 -19130 16379 -19025
rect 16476 -19029 16480 -19004
rect 16506 -19029 16510 -19004
rect 16437 -19040 16441 -19033
rect 16498 -19040 16502 -19033
rect 16430 -19043 16511 -19040
rect 16318 -19133 16379 -19130
rect 16318 -19137 16321 -19133
rect 16227 -19141 16240 -19137
rect 16236 -19160 16240 -19141
rect 16247 -19144 16251 -19137
rect 16311 -19145 16314 -19141
rect 16247 -19156 16251 -19149
rect 16304 -19148 16330 -19145
rect 16170 -19178 16174 -19164
rect 16186 -19178 16190 -19164
rect 16224 -19178 16228 -19164
rect 16244 -19178 16248 -19164
rect 16304 -19178 16307 -19148
rect 15437 -19181 16307 -19178
rect 16326 -19221 16330 -19148
rect 16617 -19156 16622 -19004
rect 16803 -19092 16809 -18971
rect 16803 -19124 16809 -19099
rect 16730 -19129 16809 -19124
rect 16736 -19141 16740 -19129
rect 16617 -19160 16737 -19156
rect 16754 -19161 16758 -19147
rect 16617 -19167 16747 -19163
rect 16754 -19165 16766 -19161
rect 15799 -19249 16081 -19244
rect 16130 -19273 16309 -19269
rect 16130 -19280 16134 -19273
rect 15853 -19283 16134 -19280
rect 15854 -19288 15859 -19283
rect 15673 -19292 15859 -19288
rect 15673 -19294 15677 -19292
rect 15501 -19297 15677 -19294
rect 15507 -19312 15511 -19297
rect 15526 -19312 15530 -19297
rect 15400 -19320 15496 -19316
rect 15550 -19312 15554 -19297
rect 15709 -19307 15713 -19292
rect 15728 -19307 15732 -19292
rect 15762 -19307 15766 -19292
rect 15964 -19298 15968 -19283
rect 15983 -19298 15987 -19283
rect 16003 -19298 16007 -19283
rect 16025 -19298 16029 -19283
rect 16225 -19288 16229 -19273
rect 16244 -19288 16248 -19273
rect 16264 -19288 16268 -19273
rect 16298 -19288 16302 -19273
rect 15633 -19311 15692 -19308
rect 15492 -19326 15496 -19320
rect 15516 -19326 15520 -19318
rect 15558 -19326 15562 -19318
rect 15688 -19321 15692 -19311
rect 15718 -19321 15722 -19313
rect 15738 -19321 15742 -19313
rect 15770 -19321 15774 -19313
rect 15973 -19312 15977 -19304
rect 15993 -19312 15997 -19304
rect 16033 -19312 16037 -19304
rect 16234 -19302 16238 -19294
rect 16254 -19302 16258 -19294
rect 16274 -19302 16278 -19294
rect 16306 -19302 16310 -19294
rect 16087 -19306 16226 -19302
rect 16234 -19306 16299 -19302
rect 16306 -19306 16357 -19302
rect 15906 -19316 15965 -19312
rect 15973 -19316 16026 -19312
rect 16033 -19316 16059 -19312
rect 15688 -19325 15710 -19321
rect 15718 -19325 15763 -19321
rect 15770 -19325 15827 -19321
rect 15492 -19330 15508 -19326
rect 15516 -19330 15551 -19326
rect 15558 -19330 15578 -19326
rect 15475 -19339 15518 -19335
rect 15526 -19344 15530 -19330
rect 15558 -19344 15562 -19330
rect 15655 -19332 15720 -19328
rect 15668 -19337 15730 -19335
rect 15673 -19339 15730 -19337
rect 15738 -19342 15742 -19325
rect 15770 -19342 15774 -19325
rect 15923 -19323 15975 -19319
rect 15930 -19330 15985 -19326
rect 15930 -19335 15934 -19330
rect 15858 -19338 15934 -19335
rect 15953 -19337 15995 -19333
rect 15953 -19342 15957 -19337
rect 16003 -19341 16007 -19316
rect 16033 -19341 16037 -19316
rect 16116 -19313 16236 -19309
rect 16133 -19320 16246 -19316
rect 16148 -19327 16256 -19323
rect 16148 -19328 16211 -19327
rect 16214 -19335 16266 -19331
rect 16214 -19337 16219 -19335
rect 15507 -19355 15511 -19348
rect 15550 -19355 15554 -19348
rect 15709 -19353 15713 -19346
rect 15762 -19353 15766 -19346
rect 15927 -19346 15957 -19342
rect 16274 -19338 16278 -19306
rect 16306 -19338 16310 -19306
rect 15964 -19352 15968 -19345
rect 16025 -19352 16029 -19345
rect 16225 -19349 16229 -19342
rect 16298 -19349 16302 -19342
rect 16552 -19343 16557 -19273
rect 16480 -19347 16557 -19343
rect 16130 -19352 16312 -19349
rect 15930 -19353 16312 -19352
rect 15700 -19355 16134 -19353
rect 15494 -19356 16134 -19355
rect 15494 -19357 15945 -19356
rect 15494 -19358 15711 -19357
rect 16486 -19359 16490 -19347
rect 16534 -19359 16538 -19347
rect 15584 -19374 15969 -19372
rect 15584 -19378 16487 -19374
rect 16524 -19379 16528 -19365
rect 16542 -19379 16546 -19365
rect 16617 -19379 16622 -19167
rect 16754 -19171 16758 -19165
rect 16745 -19175 16758 -19171
rect 16745 -19179 16749 -19175
rect 16736 -19190 16740 -19183
rect 16754 -19190 16758 -19183
rect 16729 -19194 16762 -19190
rect 15833 -19385 16497 -19381
rect 16524 -19383 16535 -19379
rect 16542 -19383 16622 -19379
rect 16803 -19268 16809 -19129
rect 16873 -19189 16879 -19045
rect 16873 -19221 16879 -19194
rect 16066 -19392 16507 -19388
rect 16364 -19399 16516 -19395
rect 16524 -19403 16528 -19383
rect 16495 -19407 16528 -19403
rect 16495 -19411 16499 -19407
rect 16514 -19411 16518 -19407
rect 16542 -19411 16546 -19383
rect 16486 -19422 16490 -19415
rect 16504 -19422 16508 -19415
rect 16524 -19422 16528 -19415
rect 16534 -19422 16538 -19415
rect 16319 -19426 16557 -19422
rect 16803 -19466 16809 -19274
rect 15551 -19469 16810 -19466
rect 15568 -19475 15571 -19469
rect 15624 -19475 15627 -19469
rect 15821 -19475 15824 -19469
rect 16084 -19475 16087 -19469
rect 15356 -19490 15564 -19487
rect 15358 -19491 15564 -19490
rect 15575 -19488 15578 -19479
rect 15575 -19491 15582 -19488
rect 15575 -19495 15578 -19491
rect 15611 -19491 15620 -19487
rect 15631 -19488 15634 -19479
rect 15631 -19491 15648 -19488
rect 15797 -19491 15817 -19487
rect 15828 -19488 15831 -19479
rect 15828 -19491 15853 -19488
rect 15631 -19495 15634 -19491
rect 15828 -19495 15831 -19491
rect 16055 -19491 16080 -19487
rect 16091 -19488 16094 -19479
rect 16091 -19491 16190 -19488
rect 16091 -19495 16094 -19491
rect 15568 -19503 15571 -19499
rect 15624 -19503 15627 -19499
rect 15821 -19503 15824 -19499
rect 16084 -19503 16087 -19499
rect 16873 -19503 16879 -19227
rect 15561 -19506 16312 -19503
rect 15582 -19507 15586 -19506
rect 16319 -19506 16879 -19503
<< m2contact >>
rect 15627 -19005 15634 -19000
rect 15876 -19012 15882 -19007
rect 16120 -19020 16127 -19014
rect 16303 -19099 16308 -19094
rect 15477 -19133 15482 -19128
rect 15436 -19149 15441 -19144
rect 15538 -19133 15543 -19128
rect 15627 -19134 15632 -19129
rect 15726 -19133 15731 -19128
rect 15518 -19149 15523 -19144
rect 15685 -19149 15690 -19144
rect 15787 -19133 15792 -19128
rect 15876 -19134 15881 -19129
rect 15983 -19133 15988 -19128
rect 15767 -19149 15772 -19144
rect 15942 -19149 15947 -19144
rect 16044 -19133 16049 -19128
rect 16120 -19134 16125 -19129
rect 16205 -19133 16210 -19128
rect 16024 -19149 16029 -19144
rect 16140 -19142 16146 -19137
rect 16154 -19150 16160 -19145
rect 16164 -19149 16169 -19144
rect 16266 -19133 16271 -19128
rect 16511 -19044 16517 -19039
rect 16246 -19149 16251 -19144
rect 16802 -19099 16809 -19092
rect 16324 -19226 16330 -19221
rect 15790 -19252 15799 -19241
rect 16081 -19251 16089 -19244
rect 16309 -19273 16316 -19267
rect 16551 -19273 16558 -19268
rect 15626 -19312 15633 -19306
rect 15900 -19317 15906 -19311
rect 16081 -19307 16087 -19301
rect 15469 -19340 15475 -19334
rect 15578 -19331 15583 -19326
rect 15648 -19334 15655 -19326
rect 15827 -19326 15833 -19321
rect 15915 -19326 15923 -19319
rect 15853 -19339 15858 -19334
rect 16059 -19317 16066 -19312
rect 16109 -19315 16116 -19309
rect 16127 -19321 16133 -19316
rect 16140 -19329 16148 -19323
rect 16213 -19342 16219 -19337
rect 16357 -19307 16364 -19302
rect 15578 -19378 15584 -19372
rect 16762 -19194 16767 -19189
rect 15827 -19386 15833 -19381
rect 16873 -19045 16880 -19039
rect 16873 -19194 16882 -19189
rect 16873 -19227 16880 -19221
rect 16803 -19274 16810 -19268
rect 16059 -19393 16066 -19388
rect 16357 -19400 16364 -19395
rect 15582 -19492 15587 -19487
rect 15648 -19491 15653 -19486
rect 15853 -19492 15858 -19487
rect 16049 -19491 16055 -19486
rect 16190 -19491 16195 -19486
<< metal2 >>
rect 15482 -19133 15538 -19129
rect 15627 -19129 15632 -19005
rect 15731 -19133 15787 -19129
rect 15876 -19129 15881 -19012
rect 15441 -19149 15518 -19144
rect 15627 -19241 15632 -19134
rect 15988 -19133 16044 -19129
rect 16120 -19129 16125 -19020
rect 16517 -19044 16873 -19039
rect 16308 -19099 16802 -19094
rect 16125 -19134 16133 -19130
rect 16210 -19133 16266 -19129
rect 15690 -19149 15767 -19144
rect 15876 -19220 15881 -19134
rect 15947 -19149 16024 -19144
rect 15876 -19226 16116 -19220
rect 15627 -19245 15790 -19241
rect 15627 -19306 15632 -19245
rect 15876 -19250 15881 -19226
rect 15791 -19302 15797 -19252
rect 15876 -19255 15922 -19250
rect 15791 -19306 15906 -19302
rect 15901 -19311 15906 -19306
rect 15915 -19319 15923 -19255
rect 16081 -19301 16087 -19251
rect 16109 -19309 16116 -19226
rect 15469 -19408 15475 -19340
rect 15578 -19372 15583 -19331
rect 15469 -19411 15598 -19408
rect 15595 -19488 15598 -19411
rect 15649 -19486 15653 -19334
rect 15827 -19381 15833 -19326
rect 15587 -19491 15598 -19488
rect 15853 -19487 15858 -19339
rect 16059 -19388 16066 -19317
rect 16127 -19316 16133 -19134
rect 16140 -19323 16146 -19142
rect 16169 -19149 16246 -19144
rect 16154 -19417 16160 -19150
rect 16767 -19194 16873 -19189
rect 16330 -19226 16873 -19221
rect 16316 -19273 16551 -19269
rect 16558 -19273 16803 -19269
rect 16190 -19342 16213 -19337
rect 16154 -19422 16161 -19417
rect 16049 -19428 16161 -19422
rect 16049 -19486 16055 -19428
rect 16190 -19486 16195 -19342
rect 16357 -19395 16364 -19307
<< m123contact >>
rect 15423 -19086 15433 -19077
rect 15423 -19151 15429 -19145
rect 15645 -19142 15650 -19137
rect 15654 -19151 15660 -19145
rect 15920 -19142 15926 -19137
rect 15895 -19149 15902 -19144
rect 15668 -19342 15673 -19337
rect 15606 -19492 15611 -19487
rect 15792 -19491 15797 -19486
rect 15920 -19347 15927 -19342
rect 16312 -19354 16319 -19349
rect 16312 -19428 16319 -19422
rect 16312 -19508 16319 -19503
<< metal3 >>
rect 15606 -19081 15660 -19076
rect 15423 -19145 15429 -19086
rect 15606 -19487 15611 -19081
rect 15645 -19264 15649 -19142
rect 15654 -19145 15660 -19081
rect 15645 -19268 15673 -19264
rect 15668 -19337 15673 -19268
rect 15896 -19345 15901 -19149
rect 15792 -19349 15901 -19345
rect 15920 -19342 15926 -19142
rect 15792 -19486 15797 -19349
rect 16312 -19422 16319 -19354
rect 16312 -19503 16319 -19428
<< labels >>
rlabel metal1 15598 -19133 15601 -19130 1 n3
rlabel metal1 15436 -19099 15526 -19095 5 VDD
rlabel metal1 15576 -19111 15601 -19108 1 VDD
rlabel metal1 15576 -19148 15601 -19145 1 GND
rlabel metal1 15437 -19181 15579 -19178 1 GND
rlabel metal1 15685 -19099 15775 -19095 5 VDD
rlabel metal1 15847 -19133 15850 -19130 1 n2
rlabel metal1 15825 -19148 15850 -19145 1 GND
rlabel metal1 15825 -19111 15850 -19108 1 VDD
rlabel metal1 15686 -19181 15828 -19178 1 GND
rlabel metal1 15942 -19099 16032 -19095 5 VDD
rlabel metal1 16104 -19133 16107 -19130 7 n1
rlabel metal1 16082 -19111 16107 -19108 1 VDD
rlabel metal1 16082 -19148 16107 -19145 1 GND
rlabel metal1 15943 -19181 16085 -19178 1 GND
rlabel metal1 16326 -19133 16329 -19130 7 n0
rlabel metal1 16164 -19099 16254 -19095 5 VDD
rlabel metal1 16304 -19111 16329 -19108 1 VDD
rlabel metal1 16304 -19148 16329 -19145 1 GND
rlabel metal1 15561 -19506 15586 -19503 1 GND
rlabel metal1 15561 -19469 15586 -19466 5 VDD
rlabel metal1 15617 -19506 15642 -19503 1 GND
rlabel metal1 15617 -19469 15642 -19466 5 VDD
rlabel metal1 15814 -19506 15839 -19503 1 GND
rlabel metal1 15814 -19469 15839 -19466 5 VDD
rlabel metal1 16077 -19506 16102 -19503 1 GND
rlabel metal1 16077 -19469 16102 -19466 5 VDD
rlabel metal1 16431 -18971 16516 -18967 5 VDD
rlabel metal1 16426 -19004 16430 -19000 1 n3
rlabel metal1 16426 -19011 16430 -19007 1 n2
rlabel metal1 16426 -19018 16430 -19014 1 n1
rlabel metal1 16426 -19025 16430 -19021 1 n0
rlabel metal1 16515 -19004 16519 -19000 1 AEB
rlabel metal1 16480 -19347 16557 -19343 5 VDD
rlabel metal1 16479 -19426 16557 -19422 1 GND
rlabel metal1 16477 -19378 16481 -19374 1 y3
rlabel metal1 16477 -19385 16481 -19381 1 y2
rlabel metal1 16477 -19392 16481 -19388 1 y1
rlabel metal1 16477 -19399 16481 -19395 1 y0
rlabel metal1 16558 -19383 16562 -19379 7 AGB
rlabel metal1 16762 -19165 16766 -19161 7 ALB
rlabel metal1 16727 -19160 16731 -19156 1 AEB
rlabel metal1 16727 -19167 16731 -19163 1 AGB
rlabel metal1 16730 -19129 16764 -19124 1 VDD
rlabel metal1 16315 -19306 16320 -19302 7 y0
rlabel metal1 16214 -19306 16219 -19302 1 n3
rlabel metal1 16214 -19313 16219 -19309 1 n2
rlabel metal1 16214 -19320 16219 -19316 1 n1
rlabel metal1 15777 -19325 15782 -19321 7 y2
rlabel metal1 15698 -19325 15703 -19321 1 n3
rlabel metal1 15702 -19357 15781 -19353 1 GND
rlabel metal1 15703 -19292 15780 -19288 5 VDD
rlabel metal1 15568 -19330 15572 -19326 7 y3
rlabel metal1 15500 -19358 15569 -19355 1 GND
rlabel metal1 15501 -19297 15568 -19294 5 VDD
rlabel metal1 15958 -19283 16043 -19280 1 VDD
rlabel metal1 16043 -19316 16047 -19312 7 y1
rlabel metal1 15953 -19323 15957 -19319 1 n2
rlabel metal1 15953 -19316 15957 -19312 1 n3
rlabel metal1 15957 -19356 16044 -19352 1 GND
rlabel metal1 15496 -19330 15500 -19326 1 CompA3
rlabel metal1 15496 -19339 15500 -19335 1 CompB3not
rlabel metal1 15698 -19332 15703 -19328 1 CompB2not
rlabel metal1 15698 -19339 15703 -19335 1 CompA2
rlabel metal1 15953 -19337 15957 -19333 1 CompA1
rlabel metal1 15953 -19330 15957 -19326 1 CompB1not
rlabel metal1 16214 -19335 16219 -19331 1 CompB0not
rlabel metal1 16214 -19327 16219 -19323 1 CompA0
rlabel metal1 16206 -19273 16303 -19269 1 VDD
rlabel metal1 15430 -19141 15434 -19137 1 CompA3
rlabel metal1 15431 -19149 15435 -19145 1 CompB3
rlabel metal1 15677 -19149 15681 -19145 1 CompB2
rlabel metal1 15677 -19141 15681 -19137 1 CompA2
rlabel metal1 15934 -19141 15938 -19137 1 CompA1
rlabel metal1 15934 -19149 15938 -19145 1 CompB1
rlabel metal1 16156 -19141 16160 -19137 1 CompA0
rlabel metal1 16161 -19149 16163 -19145 1 CompB0
rlabel metal1 15561 -19491 15564 -19487 1 CompB3
rlabel metal1 15578 -19491 15581 -19488 1 CompB3not
rlabel metal1 15616 -19491 15620 -19487 1 CompB2
rlabel metal1 15639 -19491 15642 -19488 1 CompB2not
rlabel metal1 15813 -19491 15817 -19487 1 CompB1
rlabel metal1 15836 -19491 15839 -19488 1 CompB1not
rlabel metal1 16076 -19491 16080 -19487 1 CompB0
rlabel metal1 16099 -19491 16102 -19488 1 CompB0not
rlabel metal1 16445 -19043 16462 -19040 1 GND
rlabel space 16802 -19068 16809 -19055 1 VDD
rlabel space 16873 -19102 16880 -19089 1 GND
<< end >>
