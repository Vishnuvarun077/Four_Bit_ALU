magic
tech scmos
timestamp 1701449928
<< nwell >>
rect 50 25 75 41
rect 106 25 131 41
rect 13 -52 50 -34
rect 56 -52 80 -34
rect 14 -137 51 -119
rect 57 -137 81 -119
rect 14 -226 51 -208
rect 57 -226 81 -208
rect 14 -309 51 -291
rect 57 -309 81 -291
<< ntransistor >>
rect 61 11 63 15
rect 117 11 119 15
rect 24 -76 26 -72
rect 34 -76 36 -72
rect 67 -76 69 -72
rect 25 -161 27 -157
rect 35 -161 37 -157
rect 68 -161 70 -157
rect 25 -250 27 -246
rect 35 -250 37 -246
rect 68 -250 70 -246
rect 25 -333 27 -329
rect 35 -333 37 -329
rect 68 -333 70 -329
<< ptransistor >>
rect 61 31 63 35
rect 117 31 119 35
rect 24 -46 26 -40
rect 34 -46 36 -40
rect 67 -46 69 -40
rect 25 -131 27 -125
rect 35 -131 37 -125
rect 68 -131 70 -125
rect 25 -220 27 -214
rect 35 -220 37 -214
rect 68 -220 70 -214
rect 25 -303 27 -297
rect 35 -303 37 -297
rect 68 -303 70 -297
<< ndiffusion >>
rect 60 11 61 15
rect 63 11 64 15
rect 116 11 117 15
rect 119 11 120 15
rect 23 -76 24 -72
rect 26 -76 34 -72
rect 36 -76 38 -72
rect 66 -76 67 -72
rect 69 -76 70 -72
rect 24 -161 25 -157
rect 27 -161 35 -157
rect 37 -161 39 -157
rect 67 -161 68 -157
rect 70 -161 71 -157
rect 24 -250 25 -246
rect 27 -250 35 -246
rect 37 -250 39 -246
rect 67 -250 68 -246
rect 70 -250 71 -246
rect 24 -333 25 -329
rect 27 -333 35 -329
rect 37 -333 39 -329
rect 67 -333 68 -329
rect 70 -333 71 -329
<< pdiffusion >>
rect 60 31 61 35
rect 63 31 64 35
rect 116 31 117 35
rect 119 31 120 35
rect 23 -46 24 -40
rect 26 -46 28 -40
rect 32 -46 34 -40
rect 36 -46 38 -40
rect 66 -46 67 -40
rect 69 -46 70 -40
rect 24 -131 25 -125
rect 27 -131 29 -125
rect 33 -131 35 -125
rect 37 -131 39 -125
rect 67 -131 68 -125
rect 70 -131 71 -125
rect 24 -220 25 -214
rect 27 -220 29 -214
rect 33 -220 35 -214
rect 37 -220 39 -214
rect 67 -220 68 -214
rect 70 -220 71 -214
rect 24 -303 25 -297
rect 27 -303 29 -297
rect 33 -303 35 -297
rect 37 -303 39 -297
rect 67 -303 68 -297
rect 70 -303 71 -297
<< ndcontact >>
rect 56 11 60 15
rect 64 11 68 15
rect 112 11 116 15
rect 120 11 124 15
rect 19 -76 23 -72
rect 38 -76 42 -72
rect 62 -76 66 -72
rect 70 -76 74 -72
rect 20 -161 24 -157
rect 39 -161 43 -157
rect 63 -161 67 -157
rect 71 -161 75 -157
rect 20 -250 24 -246
rect 39 -250 43 -246
rect 63 -250 67 -246
rect 71 -250 75 -246
rect 20 -333 24 -329
rect 39 -333 43 -329
rect 63 -333 67 -329
rect 71 -333 75 -329
<< pdcontact >>
rect 56 31 60 35
rect 64 31 68 35
rect 112 31 116 35
rect 120 31 124 35
rect 19 -46 23 -40
rect 28 -46 32 -40
rect 38 -46 42 -40
rect 62 -46 66 -40
rect 70 -46 74 -40
rect 20 -131 24 -125
rect 29 -131 33 -125
rect 39 -131 43 -125
rect 63 -131 67 -125
rect 71 -131 75 -125
rect 20 -220 24 -214
rect 29 -220 33 -214
rect 39 -220 43 -214
rect 63 -220 67 -214
rect 71 -220 75 -214
rect 20 -303 24 -297
rect 29 -303 33 -297
rect 39 -303 43 -297
rect 63 -303 67 -297
rect 71 -303 75 -297
<< polysilicon >>
rect 61 35 63 38
rect 117 35 119 38
rect 61 22 63 31
rect 57 20 63 22
rect 61 15 63 20
rect 117 22 119 31
rect 113 20 119 22
rect 117 15 119 20
rect 61 8 63 11
rect 117 8 119 11
rect 24 -40 26 -31
rect 34 -40 36 -31
rect 67 -40 69 -31
rect 24 -72 26 -46
rect 34 -72 36 -46
rect 67 -72 69 -46
rect 24 -79 26 -76
rect 34 -79 36 -76
rect 67 -79 69 -76
rect 25 -125 27 -116
rect 35 -125 37 -116
rect 68 -125 70 -116
rect 25 -157 27 -131
rect 35 -157 37 -131
rect 68 -157 70 -131
rect 25 -164 27 -161
rect 35 -164 37 -161
rect 68 -164 70 -161
rect 25 -214 27 -205
rect 35 -214 37 -205
rect 68 -214 70 -205
rect 25 -246 27 -220
rect 35 -246 37 -220
rect 68 -246 70 -220
rect 25 -253 27 -250
rect 35 -253 37 -250
rect 68 -253 70 -250
rect 25 -297 27 -288
rect 35 -297 37 -288
rect 68 -297 70 -288
rect 25 -329 27 -303
rect 35 -329 37 -303
rect 68 -329 70 -303
rect 25 -336 27 -333
rect 35 -336 37 -333
rect 68 -336 70 -333
<< polycontact >>
rect 53 19 57 23
rect 109 19 113 23
rect 20 -58 24 -54
rect 30 -67 34 -63
rect 63 -58 67 -54
rect 21 -143 25 -139
rect 31 -152 35 -148
rect 64 -143 68 -139
rect 21 -232 25 -228
rect 31 -241 35 -237
rect 64 -232 68 -228
rect 21 -315 25 -311
rect 31 -324 35 -320
rect 64 -315 68 -311
<< metal1 >>
rect 50 41 156 44
rect 57 35 60 41
rect 113 35 116 41
rect -37 19 53 23
rect 64 22 67 31
rect 64 19 71 22
rect -37 -139 -33 19
rect 64 15 67 19
rect 103 19 109 23
rect 120 22 123 31
rect 120 19 135 22
rect 120 15 123 19
rect 57 7 60 11
rect 113 7 116 11
rect 50 4 127 7
rect 13 -25 156 -22
rect 19 -40 23 -25
rect 38 -40 42 -25
rect 62 -40 66 -25
rect 28 -54 32 -46
rect 70 -54 74 -46
rect -24 -58 20 -54
rect 28 -58 63 -54
rect 70 -58 84 -54
rect 1 -67 30 -63
rect 38 -72 42 -58
rect 70 -72 74 -58
rect 19 -83 23 -76
rect 62 -83 66 -76
rect 12 -86 127 -83
rect 127 -107 132 -106
rect 14 -110 156 -107
rect 20 -125 24 -110
rect 39 -125 43 -110
rect 63 -125 67 -110
rect 127 -111 132 -110
rect 29 -139 33 -131
rect 71 -139 75 -131
rect -37 -143 21 -139
rect 29 -143 64 -139
rect 71 -143 85 -139
rect -37 -311 -33 -143
rect 1 -152 31 -148
rect 39 -157 43 -143
rect 71 -157 75 -143
rect 20 -168 24 -161
rect 63 -168 67 -161
rect 13 -171 127 -168
rect 14 -199 156 -196
rect 20 -214 24 -199
rect 39 -214 43 -199
rect 63 -214 67 -199
rect 29 -228 33 -220
rect 71 -228 75 -220
rect -24 -232 21 -228
rect 29 -232 64 -228
rect 71 -232 85 -228
rect -12 -241 31 -237
rect 39 -246 43 -232
rect 71 -246 75 -232
rect 20 -257 24 -250
rect 63 -257 67 -250
rect 13 -260 127 -257
rect 14 -282 156 -279
rect 20 -297 24 -282
rect 39 -297 43 -282
rect 63 -297 67 -282
rect 29 -311 33 -303
rect 71 -311 75 -303
rect -37 -315 21 -311
rect 29 -315 64 -311
rect 71 -315 85 -311
rect -12 -324 31 -320
rect 39 -329 43 -315
rect 71 -329 75 -315
rect 20 -340 24 -333
rect 63 -340 67 -333
rect 13 -343 127 -340
<< m2contact >>
rect 156 41 161 46
rect 71 18 76 23
rect 98 18 103 24
rect 127 1 132 7
rect 156 -25 161 -20
rect -29 -58 -24 -53
rect 127 -87 132 -82
rect 156 -110 161 -105
rect 127 -172 132 -167
rect 156 -199 161 -194
rect -29 -232 -24 -227
rect -17 -241 -12 -236
rect 127 -261 132 -256
rect 156 -282 162 -277
rect -17 -324 -12 -319
rect 127 -343 132 -338
<< metal2 >>
rect 73 -1 76 18
rect -31 -4 76 -1
rect -29 -53 -25 -4
rect 99 -9 102 18
rect -17 -12 102 -9
rect -29 -227 -25 -58
rect -17 -236 -13 -12
rect 127 -82 132 1
rect 127 -167 132 -87
rect -17 -319 -13 -241
rect 127 -256 132 -172
rect 127 -338 132 -261
rect 156 -20 161 41
rect 156 -105 161 -25
rect 156 -194 161 -110
rect 156 -277 161 -199
<< m123contact >>
rect 135 18 140 23
rect -4 -67 1 -62
rect -4 -152 1 -147
<< metal3 >>
rect 136 -14 140 18
rect -4 -17 140 -14
rect -4 -62 1 -17
rect -4 -147 1 -67
<< labels >>
rlabel metal1 105 19 109 23 1 S1
rlabel metal1 49 19 53 23 3 S0
rlabel metal1 50 41 131 44 5 VDD
rlabel metal1 13 -25 80 -22 1 VDD
rlabel metal1 14 -110 81 -107 1 VDD
rlabel metal1 14 -199 81 -196 1 VDD
rlabel metal1 13 -171 82 -168 1 GND
rlabel metal1 13 -260 82 -257 1 GND
rlabel metal1 79 -58 84 -54 1 D0
rlabel metal1 80 -143 85 -139 1 D1
rlabel metal1 13 -343 82 -340 1 GND
rlabel metal1 14 -282 81 -279 1 VDD
rlabel metal1 80 -232 85 -228 1 D2
rlabel metal1 80 -315 85 -311 1 D3
rlabel metal1 12 -86 81 -83 1 GND
rlabel metal1 67 4 71 7 1 GND
rlabel metal1 8 -58 13 -54 3 S0not
rlabel metal1 9 -315 14 -311 3 S0
rlabel metal1 9 -324 14 -320 3 S1
rlabel metal1 9 -241 14 -237 3 S1
rlabel metal1 9 -232 14 -228 3 S0not
rlabel metal1 9 -152 14 -148 3 S1not
rlabel metal1 9 -143 14 -139 3 S0
rlabel metal1 8 -67 13 -63 3 S1not
rlabel metal1 129 19 132 22 1 S1not
<< end >>
