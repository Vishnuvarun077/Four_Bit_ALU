magic
tech scmos
timestamp 1699811320
<< nwell >>
rect 6 148 43 166
rect 49 148 73 166
rect 92 148 129 166
rect 135 148 159 166
rect 182 148 219 166
rect 225 148 249 166
rect 277 148 314 166
rect 320 148 344 166
<< ntransistor >>
rect 17 124 19 128
rect 27 124 29 128
rect 60 124 62 128
rect 103 124 105 128
rect 113 124 115 128
rect 146 124 148 128
rect 193 124 195 128
rect 203 124 205 128
rect 236 124 238 128
rect 288 124 290 128
rect 298 124 300 128
rect 331 124 333 128
<< ptransistor >>
rect 17 154 19 160
rect 27 154 29 160
rect 60 154 62 160
rect 103 154 105 160
rect 113 154 115 160
rect 146 154 148 160
rect 193 154 195 160
rect 203 154 205 160
rect 236 154 238 160
rect 288 154 290 160
rect 298 154 300 160
rect 331 154 333 160
<< ndiffusion >>
rect 16 124 17 128
rect 19 124 27 128
rect 29 124 31 128
rect 59 124 60 128
rect 62 124 63 128
rect 102 124 103 128
rect 105 124 113 128
rect 115 124 117 128
rect 145 124 146 128
rect 148 124 149 128
rect 192 124 193 128
rect 195 124 203 128
rect 205 124 207 128
rect 235 124 236 128
rect 238 124 239 128
rect 287 124 288 128
rect 290 124 298 128
rect 300 124 302 128
rect 330 124 331 128
rect 333 124 334 128
<< pdiffusion >>
rect 16 154 17 160
rect 19 154 21 160
rect 25 154 27 160
rect 29 154 31 160
rect 59 154 60 160
rect 62 154 63 160
rect 102 154 103 160
rect 105 154 107 160
rect 111 154 113 160
rect 115 154 117 160
rect 145 154 146 160
rect 148 154 149 160
rect 192 154 193 160
rect 195 154 197 160
rect 201 154 203 160
rect 205 154 207 160
rect 235 154 236 160
rect 238 154 239 160
rect 287 154 288 160
rect 290 154 292 160
rect 296 154 298 160
rect 300 154 302 160
rect 330 154 331 160
rect 333 154 334 160
<< ndcontact >>
rect 12 124 16 128
rect 31 124 35 128
rect 55 124 59 128
rect 63 124 67 128
rect 98 124 102 128
rect 117 124 121 128
rect 141 124 145 128
rect 149 124 153 128
rect 188 124 192 128
rect 207 124 211 128
rect 231 124 235 128
rect 239 124 243 128
rect 283 124 287 128
rect 302 124 306 128
rect 326 124 330 128
rect 334 124 338 128
<< pdcontact >>
rect 12 154 16 160
rect 21 154 25 160
rect 31 154 35 160
rect 55 154 59 160
rect 63 154 67 160
rect 98 154 102 160
rect 107 154 111 160
rect 117 154 121 160
rect 141 154 145 160
rect 149 154 153 160
rect 188 154 192 160
rect 197 154 201 160
rect 207 154 211 160
rect 231 154 235 160
rect 239 154 243 160
rect 283 154 287 160
rect 292 154 296 160
rect 302 154 306 160
rect 326 154 330 160
rect 334 154 338 160
<< polysilicon >>
rect 17 160 19 169
rect 27 160 29 169
rect 60 160 62 169
rect 103 160 105 169
rect 113 160 115 169
rect 146 160 148 169
rect 193 160 195 169
rect 203 160 205 169
rect 236 160 238 169
rect 288 160 290 169
rect 298 160 300 169
rect 331 160 333 169
rect 17 128 19 154
rect 27 128 29 154
rect 60 128 62 154
rect 103 128 105 154
rect 113 128 115 154
rect 146 128 148 154
rect 193 128 195 154
rect 203 128 205 154
rect 236 128 238 154
rect 288 128 290 154
rect 298 128 300 154
rect 331 128 333 154
rect 17 121 19 124
rect 27 121 29 124
rect 60 121 62 124
rect 103 121 105 124
rect 113 121 115 124
rect 146 121 148 124
rect 193 121 195 124
rect 203 121 205 124
rect 236 121 238 124
rect 288 121 290 124
rect 298 121 300 124
rect 331 121 333 124
<< polycontact >>
rect 13 142 17 146
rect 23 133 27 137
rect 56 142 60 146
rect 99 142 103 146
rect 109 133 113 137
rect 142 142 146 146
rect 189 142 193 146
rect 199 133 203 137
rect 232 142 236 146
rect 284 142 288 146
rect 294 133 298 137
rect 327 142 331 146
<< metal1 >>
rect 6 175 344 178
rect 12 160 16 175
rect 31 160 35 175
rect 55 160 59 175
rect 98 160 102 175
rect 117 160 121 175
rect 141 160 145 175
rect 188 160 192 175
rect 207 160 211 175
rect 231 160 235 175
rect 283 160 287 175
rect 302 160 306 175
rect 326 160 330 175
rect 21 146 25 154
rect 63 146 67 154
rect 107 146 111 154
rect 149 146 153 154
rect 197 146 201 154
rect 239 146 243 154
rect 292 146 296 154
rect 334 146 338 154
rect 1 142 13 146
rect 21 142 56 146
rect 63 142 76 146
rect 87 142 99 146
rect 107 142 142 146
rect 149 142 162 146
rect 177 142 189 146
rect 197 142 232 146
rect 239 142 252 146
rect 272 142 284 146
rect 292 142 327 146
rect 334 142 347 146
rect 1 133 23 137
rect 31 128 35 142
rect 63 128 67 142
rect 87 133 109 137
rect 117 128 121 142
rect 149 128 153 142
rect 177 133 199 137
rect 207 128 211 142
rect 239 128 243 142
rect 272 133 294 137
rect 302 128 306 142
rect 334 128 338 142
rect 12 117 16 124
rect 55 117 59 124
rect 98 117 102 124
rect 141 117 145 124
rect 188 117 192 124
rect 231 117 235 124
rect 283 117 287 124
rect 326 117 330 124
rect 5 114 345 117
<< labels >>
rlabel metal1 1 142 5 146 3 A0
rlabel metal1 1 133 5 137 3 B0
rlabel metal1 72 142 76 146 1 Y0
rlabel metal1 87 142 91 146 1 A1
rlabel metal1 87 133 91 137 1 B1
rlabel metal1 158 142 162 146 1 Y1
rlabel metal1 177 142 181 146 1 A2
rlabel metal1 177 133 181 137 1 B2
rlabel metal1 248 142 252 146 1 Y2
rlabel metal1 272 142 276 146 1 A3
rlabel metal1 272 133 276 137 1 B3
rlabel metal1 343 142 347 146 7 Y3
rlabel metal1 308 142 312 146 1 Y3not
rlabel metal1 215 142 219 146 1 Y2not
rlabel metal1 131 142 135 146 1 Y1not
rlabel metal1 45 142 49 146 1 Y0not
rlabel metal1 24 114 34 117 1 GND
rlabel metal1 98 114 108 117 1 GND
rlabel metal1 181 114 191 117 1 GND
rlabel metal1 279 114 289 117 1 GND
rlabel metal1 28 175 38 178 5 VDD
rlabel metal1 96 175 106 178 5 VDD
rlabel metal1 193 175 203 178 5 VDD
rlabel metal1 291 175 301 178 5 VDD
<< end >>
