magic
tech scmos
timestamp 1701524471
<< nwell >>
rect 1605 3390 1695 3408
rect 1767 3399 1857 3417
rect 2004 3409 2094 3427
rect 1893 3283 1930 3301
rect 1936 3283 1960 3301
rect 2021 3284 2058 3302
rect 2064 3284 2088 3302
rect 2062 3212 2119 3230
rect 1614 3058 1704 3076
rect 1776 3067 1866 3085
rect 2013 3077 2103 3095
rect 1902 2951 1939 2969
rect 1945 2951 1969 2969
rect 2030 2952 2067 2970
rect 2073 2952 2097 2970
rect 2071 2880 2128 2898
rect 1635 2692 1725 2710
rect 1797 2701 1887 2719
rect 2034 2711 2124 2729
rect 1923 2585 1960 2603
rect 1966 2585 1990 2603
rect 2051 2586 2088 2604
rect 2094 2586 2118 2604
rect 2092 2514 2149 2532
rect 1663 2318 1753 2336
rect 1825 2327 1915 2345
rect 2062 2337 2152 2355
rect 1951 2211 1988 2229
rect 1994 2211 2018 2229
rect 2079 2212 2116 2230
rect 2122 2212 2146 2230
rect 2120 2140 2177 2158
rect 3948 1775 4003 1793
rect 4009 1775 4033 1793
rect 1042 1717 1067 1733
rect 1098 1717 1123 1733
rect 1738 1701 1775 1719
rect 1781 1701 1805 1719
rect 1824 1701 1861 1719
rect 1867 1701 1891 1719
rect 1914 1701 1951 1719
rect 1957 1701 1981 1719
rect 2009 1701 2046 1719
rect 2052 1701 2076 1719
rect 2093 1701 2130 1719
rect 2136 1701 2160 1719
rect 2179 1701 2216 1719
rect 2222 1701 2246 1719
rect 2269 1701 2306 1719
rect 2312 1701 2336 1719
rect 2364 1701 2401 1719
rect 2407 1701 2431 1719
rect 1005 1640 1042 1658
rect 1048 1640 1072 1658
rect 2953 1649 3043 1667
rect 3093 1646 3118 1662
rect 3202 1649 3292 1667
rect 3342 1646 3367 1662
rect 3459 1649 3549 1667
rect 3599 1646 3624 1662
rect 3681 1649 3771 1667
rect 3821 1646 3846 1662
rect 4247 1620 4281 1638
rect 1006 1555 1043 1573
rect 1049 1555 1073 1573
rect 1311 1569 1368 1587
rect 1006 1466 1043 1484
rect 1049 1466 1073 1484
rect 1716 1457 1753 1475
rect 1759 1457 1783 1475
rect 1802 1457 1839 1475
rect 1845 1457 1869 1475
rect 1892 1457 1929 1475
rect 1935 1457 1959 1475
rect 1987 1457 2024 1475
rect 2030 1457 2054 1475
rect 2071 1457 2108 1475
rect 2114 1457 2138 1475
rect 2157 1457 2194 1475
rect 2200 1457 2224 1475
rect 2247 1457 2284 1475
rect 2290 1457 2314 1475
rect 2342 1457 2379 1475
rect 2385 1457 2409 1475
rect 3018 1449 3055 1467
rect 3061 1449 3085 1467
rect 3220 1454 3266 1472
rect 3273 1454 3297 1472
rect 3475 1463 3530 1481
rect 3536 1463 3560 1481
rect 3736 1473 3801 1491
rect 3809 1473 3833 1491
rect 3997 1402 4074 1420
rect 1006 1383 1043 1401
rect 1049 1383 1073 1401
rect 3078 1288 3103 1304
rect 3134 1288 3159 1304
rect 3331 1288 3356 1304
rect 3594 1288 3619 1304
rect 1760 1140 1797 1158
rect 1803 1140 1827 1158
rect 1846 1140 1883 1158
rect 1889 1140 1913 1158
rect 1936 1140 1973 1158
rect 1979 1140 2003 1158
rect 2031 1140 2068 1158
rect 2074 1140 2098 1158
rect 2115 1140 2152 1158
rect 2158 1140 2182 1158
rect 2201 1140 2238 1158
rect 2244 1140 2268 1158
rect 2291 1140 2328 1158
rect 2334 1140 2358 1158
rect 2386 1140 2423 1158
rect 2429 1140 2453 1158
rect 1822 1039 1859 1057
rect 1865 1039 1889 1057
rect 1908 1039 1945 1057
rect 1951 1039 1975 1057
rect 1998 1039 2035 1057
rect 2041 1039 2065 1057
rect 2093 1039 2130 1057
rect 2136 1039 2160 1057
<< ntransistor >>
rect 1616 3350 1618 3354
rect 1632 3350 1634 3354
rect 1642 3350 1644 3354
rect 1652 3350 1654 3354
rect 1662 3350 1664 3354
rect 1778 3359 1780 3363
rect 1794 3359 1796 3363
rect 1804 3359 1806 3363
rect 1814 3359 1816 3363
rect 1824 3359 1826 3363
rect 1682 3350 1684 3354
rect 2015 3369 2017 3373
rect 2031 3369 2033 3373
rect 2041 3369 2043 3373
rect 2051 3369 2053 3373
rect 2061 3369 2063 3373
rect 1844 3359 1846 3363
rect 2081 3369 2083 3373
rect 1904 3259 1906 3263
rect 1914 3259 1916 3263
rect 1947 3259 1949 3263
rect 2032 3260 2034 3264
rect 2042 3260 2044 3264
rect 2075 3260 2077 3264
rect 2073 3182 2075 3186
rect 2083 3182 2085 3186
rect 2101 3182 2103 3186
rect 1625 3018 1627 3022
rect 1641 3018 1643 3022
rect 1651 3018 1653 3022
rect 1661 3018 1663 3022
rect 1671 3018 1673 3022
rect 1787 3027 1789 3031
rect 1803 3027 1805 3031
rect 1813 3027 1815 3031
rect 1823 3027 1825 3031
rect 1833 3027 1835 3031
rect 1691 3018 1693 3022
rect 2024 3037 2026 3041
rect 2040 3037 2042 3041
rect 2050 3037 2052 3041
rect 2060 3037 2062 3041
rect 2070 3037 2072 3041
rect 1853 3027 1855 3031
rect 2090 3037 2092 3041
rect 1913 2927 1915 2931
rect 1923 2927 1925 2931
rect 1956 2927 1958 2931
rect 2041 2928 2043 2932
rect 2051 2928 2053 2932
rect 2084 2928 2086 2932
rect 2082 2850 2084 2854
rect 2092 2850 2094 2854
rect 2110 2850 2112 2854
rect 1646 2652 1648 2656
rect 1662 2652 1664 2656
rect 1672 2652 1674 2656
rect 1682 2652 1684 2656
rect 1692 2652 1694 2656
rect 1808 2661 1810 2665
rect 1824 2661 1826 2665
rect 1834 2661 1836 2665
rect 1844 2661 1846 2665
rect 1854 2661 1856 2665
rect 1712 2652 1714 2656
rect 2045 2671 2047 2675
rect 2061 2671 2063 2675
rect 2071 2671 2073 2675
rect 2081 2671 2083 2675
rect 2091 2671 2093 2675
rect 1874 2661 1876 2665
rect 2111 2671 2113 2675
rect 1934 2561 1936 2565
rect 1944 2561 1946 2565
rect 1977 2561 1979 2565
rect 2062 2562 2064 2566
rect 2072 2562 2074 2566
rect 2105 2562 2107 2566
rect 2103 2484 2105 2488
rect 2113 2484 2115 2488
rect 2131 2484 2133 2488
rect 1674 2278 1676 2282
rect 1690 2278 1692 2282
rect 1700 2278 1702 2282
rect 1710 2278 1712 2282
rect 1720 2278 1722 2282
rect 1836 2287 1838 2291
rect 1852 2287 1854 2291
rect 1862 2287 1864 2291
rect 1872 2287 1874 2291
rect 1882 2287 1884 2291
rect 1740 2278 1742 2282
rect 2073 2297 2075 2301
rect 2089 2297 2091 2301
rect 2099 2297 2101 2301
rect 2109 2297 2111 2301
rect 2119 2297 2121 2301
rect 1902 2287 1904 2291
rect 2139 2297 2141 2301
rect 1962 2187 1964 2191
rect 1972 2187 1974 2191
rect 2005 2187 2007 2191
rect 2090 2188 2092 2192
rect 2100 2188 2102 2192
rect 2133 2188 2135 2192
rect 2131 2110 2133 2114
rect 2141 2110 2143 2114
rect 2159 2110 2161 2114
rect 3959 1740 3961 1744
rect 3969 1740 3971 1744
rect 3979 1740 3981 1744
rect 3989 1740 3991 1744
rect 4020 1740 4022 1744
rect 1053 1703 1055 1707
rect 1109 1703 1111 1707
rect 1749 1677 1751 1681
rect 1759 1677 1761 1681
rect 1792 1677 1794 1681
rect 1835 1677 1837 1681
rect 1845 1677 1847 1681
rect 1878 1677 1880 1681
rect 1925 1677 1927 1681
rect 1935 1677 1937 1681
rect 1968 1677 1970 1681
rect 2020 1677 2022 1681
rect 2030 1677 2032 1681
rect 2063 1677 2065 1681
rect 2104 1677 2106 1681
rect 2114 1677 2116 1681
rect 2147 1677 2149 1681
rect 2190 1677 2192 1681
rect 2200 1677 2202 1681
rect 2233 1677 2235 1681
rect 2280 1677 2282 1681
rect 2290 1677 2292 1681
rect 2323 1677 2325 1681
rect 2375 1677 2377 1681
rect 2385 1677 2387 1681
rect 2418 1677 2420 1681
rect 1016 1616 1018 1620
rect 1026 1616 1028 1620
rect 1059 1616 1061 1620
rect 3104 1632 3106 1636
rect 2964 1609 2966 1613
rect 2980 1609 2982 1613
rect 2990 1609 2992 1613
rect 3000 1609 3002 1613
rect 3010 1609 3012 1613
rect 3353 1632 3355 1636
rect 3030 1609 3032 1613
rect 3213 1609 3215 1613
rect 3229 1609 3231 1613
rect 3239 1609 3241 1613
rect 3249 1609 3251 1613
rect 3259 1609 3261 1613
rect 3610 1632 3612 1636
rect 3279 1609 3281 1613
rect 3470 1609 3472 1613
rect 3486 1609 3488 1613
rect 3496 1609 3498 1613
rect 3506 1609 3508 1613
rect 3516 1609 3518 1613
rect 3832 1632 3834 1636
rect 3536 1609 3538 1613
rect 3692 1609 3694 1613
rect 3708 1609 3710 1613
rect 3718 1609 3720 1613
rect 3728 1609 3730 1613
rect 3738 1609 3740 1613
rect 3758 1609 3760 1613
rect 4258 1590 4260 1594
rect 4268 1590 4270 1594
rect 1322 1539 1324 1543
rect 1332 1539 1334 1543
rect 1350 1539 1352 1543
rect 1017 1531 1019 1535
rect 1027 1531 1029 1535
rect 1060 1531 1062 1535
rect 1017 1442 1019 1446
rect 1027 1442 1029 1446
rect 1060 1442 1062 1446
rect 1727 1433 1729 1437
rect 1737 1433 1739 1437
rect 1770 1433 1772 1437
rect 1813 1433 1815 1437
rect 1823 1433 1825 1437
rect 1856 1433 1858 1437
rect 1903 1433 1905 1437
rect 1913 1433 1915 1437
rect 1946 1433 1948 1437
rect 1998 1433 2000 1437
rect 2008 1433 2010 1437
rect 2041 1433 2043 1437
rect 2082 1433 2084 1437
rect 2092 1433 2094 1437
rect 2125 1433 2127 1437
rect 2168 1433 2170 1437
rect 2178 1433 2180 1437
rect 2211 1433 2213 1437
rect 2258 1433 2260 1437
rect 2268 1433 2270 1437
rect 2301 1433 2303 1437
rect 2353 1433 2355 1437
rect 2363 1433 2365 1437
rect 2396 1433 2398 1437
rect 3029 1425 3031 1429
rect 3039 1425 3041 1429
rect 3072 1425 3074 1429
rect 3231 1427 3233 1431
rect 3241 1427 3243 1431
rect 3251 1427 3253 1431
rect 3284 1427 3286 1431
rect 3486 1428 3488 1432
rect 3496 1428 3498 1432
rect 3506 1428 3508 1432
rect 3516 1428 3518 1432
rect 3547 1428 3549 1432
rect 3747 1431 3749 1435
rect 3757 1431 3759 1435
rect 3767 1431 3769 1435
rect 3777 1431 3779 1435
rect 3787 1431 3789 1435
rect 3820 1431 3822 1435
rect 1017 1359 1019 1363
rect 1027 1359 1029 1363
rect 1060 1359 1062 1363
rect 4008 1358 4010 1362
rect 4018 1358 4020 1362
rect 4027 1358 4029 1362
rect 4037 1358 4039 1362
rect 4056 1358 4058 1362
rect 3089 1274 3091 1278
rect 3145 1274 3147 1278
rect 3342 1274 3344 1278
rect 3605 1274 3607 1278
rect 1771 1116 1773 1120
rect 1781 1116 1783 1120
rect 1814 1116 1816 1120
rect 1857 1116 1859 1120
rect 1867 1116 1869 1120
rect 1900 1116 1902 1120
rect 1947 1116 1949 1120
rect 1957 1116 1959 1120
rect 1990 1116 1992 1120
rect 2042 1116 2044 1120
rect 2052 1116 2054 1120
rect 2085 1116 2087 1120
rect 2126 1116 2128 1120
rect 2136 1116 2138 1120
rect 2169 1116 2171 1120
rect 2212 1116 2214 1120
rect 2222 1116 2224 1120
rect 2255 1116 2257 1120
rect 2302 1116 2304 1120
rect 2312 1116 2314 1120
rect 2345 1116 2347 1120
rect 2397 1116 2399 1120
rect 2407 1116 2409 1120
rect 2440 1116 2442 1120
rect 1833 1015 1835 1019
rect 1843 1015 1845 1019
rect 1876 1015 1878 1019
rect 1919 1015 1921 1019
rect 1929 1015 1931 1019
rect 1962 1015 1964 1019
rect 2009 1015 2011 1019
rect 2019 1015 2021 1019
rect 2052 1015 2054 1019
rect 2104 1015 2106 1019
rect 2114 1015 2116 1019
rect 2147 1015 2149 1019
<< ptransistor >>
rect 1616 3396 1618 3402
rect 1632 3396 1634 3402
rect 1642 3396 1644 3402
rect 1652 3396 1654 3402
rect 1662 3396 1664 3402
rect 1682 3396 1684 3402
rect 1778 3405 1780 3411
rect 1794 3405 1796 3411
rect 1804 3405 1806 3411
rect 1814 3405 1816 3411
rect 1824 3405 1826 3411
rect 1844 3405 1846 3411
rect 2015 3415 2017 3421
rect 2031 3415 2033 3421
rect 2041 3415 2043 3421
rect 2051 3415 2053 3421
rect 2061 3415 2063 3421
rect 2081 3415 2083 3421
rect 1904 3289 1906 3295
rect 1914 3289 1916 3295
rect 1947 3289 1949 3295
rect 2032 3290 2034 3296
rect 2042 3290 2044 3296
rect 2075 3290 2077 3296
rect 2073 3218 2075 3224
rect 2083 3218 2085 3224
rect 2101 3218 2103 3224
rect 1625 3064 1627 3070
rect 1641 3064 1643 3070
rect 1651 3064 1653 3070
rect 1661 3064 1663 3070
rect 1671 3064 1673 3070
rect 1691 3064 1693 3070
rect 1787 3073 1789 3079
rect 1803 3073 1805 3079
rect 1813 3073 1815 3079
rect 1823 3073 1825 3079
rect 1833 3073 1835 3079
rect 1853 3073 1855 3079
rect 2024 3083 2026 3089
rect 2040 3083 2042 3089
rect 2050 3083 2052 3089
rect 2060 3083 2062 3089
rect 2070 3083 2072 3089
rect 2090 3083 2092 3089
rect 1913 2957 1915 2963
rect 1923 2957 1925 2963
rect 1956 2957 1958 2963
rect 2041 2958 2043 2964
rect 2051 2958 2053 2964
rect 2084 2958 2086 2964
rect 2082 2886 2084 2892
rect 2092 2886 2094 2892
rect 2110 2886 2112 2892
rect 1646 2698 1648 2704
rect 1662 2698 1664 2704
rect 1672 2698 1674 2704
rect 1682 2698 1684 2704
rect 1692 2698 1694 2704
rect 1712 2698 1714 2704
rect 1808 2707 1810 2713
rect 1824 2707 1826 2713
rect 1834 2707 1836 2713
rect 1844 2707 1846 2713
rect 1854 2707 1856 2713
rect 1874 2707 1876 2713
rect 2045 2717 2047 2723
rect 2061 2717 2063 2723
rect 2071 2717 2073 2723
rect 2081 2717 2083 2723
rect 2091 2717 2093 2723
rect 2111 2717 2113 2723
rect 1934 2591 1936 2597
rect 1944 2591 1946 2597
rect 1977 2591 1979 2597
rect 2062 2592 2064 2598
rect 2072 2592 2074 2598
rect 2105 2592 2107 2598
rect 2103 2520 2105 2526
rect 2113 2520 2115 2526
rect 2131 2520 2133 2526
rect 1674 2324 1676 2330
rect 1690 2324 1692 2330
rect 1700 2324 1702 2330
rect 1710 2324 1712 2330
rect 1720 2324 1722 2330
rect 1740 2324 1742 2330
rect 1836 2333 1838 2339
rect 1852 2333 1854 2339
rect 1862 2333 1864 2339
rect 1872 2333 1874 2339
rect 1882 2333 1884 2339
rect 1902 2333 1904 2339
rect 2073 2343 2075 2349
rect 2089 2343 2091 2349
rect 2099 2343 2101 2349
rect 2109 2343 2111 2349
rect 2119 2343 2121 2349
rect 2139 2343 2141 2349
rect 1962 2217 1964 2223
rect 1972 2217 1974 2223
rect 2005 2217 2007 2223
rect 2090 2218 2092 2224
rect 2100 2218 2102 2224
rect 2133 2218 2135 2224
rect 2131 2146 2133 2152
rect 2141 2146 2143 2152
rect 2159 2146 2161 2152
rect 3959 1781 3961 1787
rect 3969 1781 3971 1787
rect 3979 1781 3981 1787
rect 3989 1781 3991 1787
rect 4020 1781 4022 1787
rect 1053 1723 1055 1727
rect 1109 1723 1111 1727
rect 1749 1707 1751 1713
rect 1759 1707 1761 1713
rect 1792 1707 1794 1713
rect 1835 1707 1837 1713
rect 1845 1707 1847 1713
rect 1878 1707 1880 1713
rect 1925 1707 1927 1713
rect 1935 1707 1937 1713
rect 1968 1707 1970 1713
rect 2020 1707 2022 1713
rect 2030 1707 2032 1713
rect 2063 1707 2065 1713
rect 2104 1707 2106 1713
rect 2114 1707 2116 1713
rect 2147 1707 2149 1713
rect 2190 1707 2192 1713
rect 2200 1707 2202 1713
rect 2233 1707 2235 1713
rect 2280 1707 2282 1713
rect 2290 1707 2292 1713
rect 2323 1707 2325 1713
rect 2375 1707 2377 1713
rect 2385 1707 2387 1713
rect 2418 1707 2420 1713
rect 2964 1655 2966 1661
rect 2980 1655 2982 1661
rect 2990 1655 2992 1661
rect 3000 1655 3002 1661
rect 3010 1655 3012 1661
rect 3030 1655 3032 1661
rect 1016 1646 1018 1652
rect 1026 1646 1028 1652
rect 1059 1646 1061 1652
rect 3104 1652 3106 1656
rect 3213 1655 3215 1661
rect 3229 1655 3231 1661
rect 3239 1655 3241 1661
rect 3249 1655 3251 1661
rect 3259 1655 3261 1661
rect 3279 1655 3281 1661
rect 3353 1652 3355 1656
rect 3470 1655 3472 1661
rect 3486 1655 3488 1661
rect 3496 1655 3498 1661
rect 3506 1655 3508 1661
rect 3516 1655 3518 1661
rect 3536 1655 3538 1661
rect 3610 1652 3612 1656
rect 3692 1655 3694 1661
rect 3708 1655 3710 1661
rect 3718 1655 3720 1661
rect 3728 1655 3730 1661
rect 3738 1655 3740 1661
rect 3758 1655 3760 1661
rect 3832 1652 3834 1656
rect 4258 1626 4260 1632
rect 4268 1626 4270 1632
rect 1322 1575 1324 1581
rect 1332 1575 1334 1581
rect 1350 1575 1352 1581
rect 1017 1561 1019 1567
rect 1027 1561 1029 1567
rect 1060 1561 1062 1567
rect 1017 1472 1019 1478
rect 1027 1472 1029 1478
rect 1060 1472 1062 1478
rect 3747 1479 3749 1485
rect 3757 1479 3759 1485
rect 3767 1479 3769 1485
rect 3777 1479 3779 1485
rect 3787 1479 3789 1485
rect 3820 1479 3822 1485
rect 1727 1463 1729 1469
rect 1737 1463 1739 1469
rect 1770 1463 1772 1469
rect 1813 1463 1815 1469
rect 1823 1463 1825 1469
rect 1856 1463 1858 1469
rect 1903 1463 1905 1469
rect 1913 1463 1915 1469
rect 1946 1463 1948 1469
rect 1998 1463 2000 1469
rect 2008 1463 2010 1469
rect 2041 1463 2043 1469
rect 2082 1463 2084 1469
rect 2092 1463 2094 1469
rect 2125 1463 2127 1469
rect 2168 1463 2170 1469
rect 2178 1463 2180 1469
rect 2211 1463 2213 1469
rect 2258 1463 2260 1469
rect 2268 1463 2270 1469
rect 2301 1463 2303 1469
rect 2353 1463 2355 1469
rect 2363 1463 2365 1469
rect 2396 1463 2398 1469
rect 3486 1469 3488 1475
rect 3496 1469 3498 1475
rect 3506 1469 3508 1475
rect 3516 1469 3518 1475
rect 3547 1469 3549 1475
rect 3029 1455 3031 1461
rect 3039 1455 3041 1461
rect 3072 1455 3074 1461
rect 3231 1460 3233 1466
rect 3241 1460 3243 1466
rect 3251 1460 3253 1466
rect 3284 1460 3286 1466
rect 4008 1408 4010 1414
rect 4018 1408 4020 1414
rect 4027 1408 4029 1414
rect 4037 1408 4039 1414
rect 4056 1408 4058 1414
rect 1017 1389 1019 1395
rect 1027 1389 1029 1395
rect 1060 1389 1062 1395
rect 3089 1294 3091 1298
rect 3145 1294 3147 1298
rect 3342 1294 3344 1298
rect 3605 1294 3607 1298
rect 1771 1146 1773 1152
rect 1781 1146 1783 1152
rect 1814 1146 1816 1152
rect 1857 1146 1859 1152
rect 1867 1146 1869 1152
rect 1900 1146 1902 1152
rect 1947 1146 1949 1152
rect 1957 1146 1959 1152
rect 1990 1146 1992 1152
rect 2042 1146 2044 1152
rect 2052 1146 2054 1152
rect 2085 1146 2087 1152
rect 2126 1146 2128 1152
rect 2136 1146 2138 1152
rect 2169 1146 2171 1152
rect 2212 1146 2214 1152
rect 2222 1146 2224 1152
rect 2255 1146 2257 1152
rect 2302 1146 2304 1152
rect 2312 1146 2314 1152
rect 2345 1146 2347 1152
rect 2397 1146 2399 1152
rect 2407 1146 2409 1152
rect 2440 1146 2442 1152
rect 1833 1045 1835 1051
rect 1843 1045 1845 1051
rect 1876 1045 1878 1051
rect 1919 1045 1921 1051
rect 1929 1045 1931 1051
rect 1962 1045 1964 1051
rect 2009 1045 2011 1051
rect 2019 1045 2021 1051
rect 2052 1045 2054 1051
rect 2104 1045 2106 1051
rect 2114 1045 2116 1051
rect 2147 1045 2149 1051
<< ndiffusion >>
rect 1615 3350 1616 3354
rect 1618 3350 1619 3354
rect 1631 3350 1632 3354
rect 1634 3350 1642 3354
rect 1644 3350 1646 3354
rect 1650 3350 1652 3354
rect 1654 3350 1662 3354
rect 1664 3350 1665 3354
rect 1777 3359 1778 3363
rect 1780 3359 1781 3363
rect 1793 3359 1794 3363
rect 1796 3359 1804 3363
rect 1806 3359 1808 3363
rect 1812 3359 1814 3363
rect 1816 3359 1824 3363
rect 1826 3359 1827 3363
rect 1681 3350 1682 3354
rect 1684 3350 1685 3354
rect 2014 3369 2015 3373
rect 2017 3369 2018 3373
rect 2030 3369 2031 3373
rect 2033 3369 2041 3373
rect 2043 3369 2045 3373
rect 2049 3369 2051 3373
rect 2053 3369 2061 3373
rect 2063 3369 2064 3373
rect 1843 3359 1844 3363
rect 1846 3359 1847 3363
rect 2080 3369 2081 3373
rect 2083 3369 2084 3373
rect 1903 3259 1904 3263
rect 1906 3259 1914 3263
rect 1916 3259 1918 3263
rect 1946 3259 1947 3263
rect 1949 3259 1950 3263
rect 2031 3260 2032 3264
rect 2034 3260 2042 3264
rect 2044 3260 2046 3264
rect 2074 3260 2075 3264
rect 2077 3260 2078 3264
rect 2072 3182 2073 3186
rect 2075 3182 2077 3186
rect 2081 3182 2083 3186
rect 2085 3182 2086 3186
rect 2100 3182 2101 3186
rect 2103 3182 2104 3186
rect 1624 3018 1625 3022
rect 1627 3018 1628 3022
rect 1640 3018 1641 3022
rect 1643 3018 1651 3022
rect 1653 3018 1655 3022
rect 1659 3018 1661 3022
rect 1663 3018 1671 3022
rect 1673 3018 1674 3022
rect 1786 3027 1787 3031
rect 1789 3027 1790 3031
rect 1802 3027 1803 3031
rect 1805 3027 1813 3031
rect 1815 3027 1817 3031
rect 1821 3027 1823 3031
rect 1825 3027 1833 3031
rect 1835 3027 1836 3031
rect 1690 3018 1691 3022
rect 1693 3018 1694 3022
rect 2023 3037 2024 3041
rect 2026 3037 2027 3041
rect 2039 3037 2040 3041
rect 2042 3037 2050 3041
rect 2052 3037 2054 3041
rect 2058 3037 2060 3041
rect 2062 3037 2070 3041
rect 2072 3037 2073 3041
rect 1852 3027 1853 3031
rect 1855 3027 1856 3031
rect 2089 3037 2090 3041
rect 2092 3037 2093 3041
rect 1912 2927 1913 2931
rect 1915 2927 1923 2931
rect 1925 2927 1927 2931
rect 1955 2927 1956 2931
rect 1958 2927 1959 2931
rect 2040 2928 2041 2932
rect 2043 2928 2051 2932
rect 2053 2928 2055 2932
rect 2083 2928 2084 2932
rect 2086 2928 2087 2932
rect 2081 2850 2082 2854
rect 2084 2850 2086 2854
rect 2090 2850 2092 2854
rect 2094 2850 2095 2854
rect 2109 2850 2110 2854
rect 2112 2850 2113 2854
rect 1645 2652 1646 2656
rect 1648 2652 1649 2656
rect 1661 2652 1662 2656
rect 1664 2652 1672 2656
rect 1674 2652 1676 2656
rect 1680 2652 1682 2656
rect 1684 2652 1692 2656
rect 1694 2652 1695 2656
rect 1807 2661 1808 2665
rect 1810 2661 1811 2665
rect 1823 2661 1824 2665
rect 1826 2661 1834 2665
rect 1836 2661 1838 2665
rect 1842 2661 1844 2665
rect 1846 2661 1854 2665
rect 1856 2661 1857 2665
rect 1711 2652 1712 2656
rect 1714 2652 1715 2656
rect 2044 2671 2045 2675
rect 2047 2671 2048 2675
rect 2060 2671 2061 2675
rect 2063 2671 2071 2675
rect 2073 2671 2075 2675
rect 2079 2671 2081 2675
rect 2083 2671 2091 2675
rect 2093 2671 2094 2675
rect 1873 2661 1874 2665
rect 1876 2661 1877 2665
rect 2110 2671 2111 2675
rect 2113 2671 2114 2675
rect 1933 2561 1934 2565
rect 1936 2561 1944 2565
rect 1946 2561 1948 2565
rect 1976 2561 1977 2565
rect 1979 2561 1980 2565
rect 2061 2562 2062 2566
rect 2064 2562 2072 2566
rect 2074 2562 2076 2566
rect 2104 2562 2105 2566
rect 2107 2562 2108 2566
rect 2102 2484 2103 2488
rect 2105 2484 2107 2488
rect 2111 2484 2113 2488
rect 2115 2484 2116 2488
rect 2130 2484 2131 2488
rect 2133 2484 2134 2488
rect 1673 2278 1674 2282
rect 1676 2278 1677 2282
rect 1689 2278 1690 2282
rect 1692 2278 1700 2282
rect 1702 2278 1704 2282
rect 1708 2278 1710 2282
rect 1712 2278 1720 2282
rect 1722 2278 1723 2282
rect 1835 2287 1836 2291
rect 1838 2287 1839 2291
rect 1851 2287 1852 2291
rect 1854 2287 1862 2291
rect 1864 2287 1866 2291
rect 1870 2287 1872 2291
rect 1874 2287 1882 2291
rect 1884 2287 1885 2291
rect 1739 2278 1740 2282
rect 1742 2278 1743 2282
rect 2072 2297 2073 2301
rect 2075 2297 2076 2301
rect 2088 2297 2089 2301
rect 2091 2297 2099 2301
rect 2101 2297 2103 2301
rect 2107 2297 2109 2301
rect 2111 2297 2119 2301
rect 2121 2297 2122 2301
rect 1901 2287 1902 2291
rect 1904 2287 1905 2291
rect 2138 2297 2139 2301
rect 2141 2297 2142 2301
rect 1961 2187 1962 2191
rect 1964 2187 1972 2191
rect 1974 2187 1976 2191
rect 2004 2187 2005 2191
rect 2007 2187 2008 2191
rect 2089 2188 2090 2192
rect 2092 2188 2100 2192
rect 2102 2188 2104 2192
rect 2132 2188 2133 2192
rect 2135 2188 2136 2192
rect 2130 2110 2131 2114
rect 2133 2110 2135 2114
rect 2139 2110 2141 2114
rect 2143 2110 2144 2114
rect 2158 2110 2159 2114
rect 2161 2110 2162 2114
rect 3958 1740 3959 1744
rect 3961 1740 3969 1744
rect 3971 1740 3979 1744
rect 3981 1740 3989 1744
rect 3991 1740 3993 1744
rect 4019 1740 4020 1744
rect 4022 1740 4023 1744
rect 1052 1703 1053 1707
rect 1055 1703 1056 1707
rect 1108 1703 1109 1707
rect 1111 1703 1112 1707
rect 1748 1677 1749 1681
rect 1751 1677 1759 1681
rect 1761 1677 1763 1681
rect 1791 1677 1792 1681
rect 1794 1677 1795 1681
rect 1834 1677 1835 1681
rect 1837 1677 1845 1681
rect 1847 1677 1849 1681
rect 1877 1677 1878 1681
rect 1880 1677 1881 1681
rect 1924 1677 1925 1681
rect 1927 1677 1935 1681
rect 1937 1677 1939 1681
rect 1967 1677 1968 1681
rect 1970 1677 1971 1681
rect 2019 1677 2020 1681
rect 2022 1677 2030 1681
rect 2032 1677 2034 1681
rect 2062 1677 2063 1681
rect 2065 1677 2066 1681
rect 2103 1677 2104 1681
rect 2106 1677 2114 1681
rect 2116 1677 2118 1681
rect 2146 1677 2147 1681
rect 2149 1677 2150 1681
rect 2189 1677 2190 1681
rect 2192 1677 2200 1681
rect 2202 1677 2204 1681
rect 2232 1677 2233 1681
rect 2235 1677 2236 1681
rect 2279 1677 2280 1681
rect 2282 1677 2290 1681
rect 2292 1677 2294 1681
rect 2322 1677 2323 1681
rect 2325 1677 2326 1681
rect 2374 1677 2375 1681
rect 2377 1677 2385 1681
rect 2387 1677 2389 1681
rect 2417 1677 2418 1681
rect 2420 1677 2421 1681
rect 1015 1616 1016 1620
rect 1018 1616 1026 1620
rect 1028 1616 1030 1620
rect 1058 1616 1059 1620
rect 1061 1616 1062 1620
rect 3103 1632 3104 1636
rect 3106 1632 3107 1636
rect 2963 1609 2964 1613
rect 2966 1609 2967 1613
rect 2979 1609 2980 1613
rect 2982 1609 2990 1613
rect 2992 1609 2994 1613
rect 2998 1609 3000 1613
rect 3002 1609 3010 1613
rect 3012 1609 3013 1613
rect 3352 1632 3353 1636
rect 3355 1632 3356 1636
rect 3029 1609 3030 1613
rect 3032 1609 3033 1613
rect 3212 1609 3213 1613
rect 3215 1609 3216 1613
rect 3228 1609 3229 1613
rect 3231 1609 3239 1613
rect 3241 1609 3243 1613
rect 3247 1609 3249 1613
rect 3251 1609 3259 1613
rect 3261 1609 3262 1613
rect 3609 1632 3610 1636
rect 3612 1632 3613 1636
rect 3278 1609 3279 1613
rect 3281 1609 3282 1613
rect 3469 1609 3470 1613
rect 3472 1609 3473 1613
rect 3485 1609 3486 1613
rect 3488 1609 3496 1613
rect 3498 1609 3500 1613
rect 3504 1609 3506 1613
rect 3508 1609 3516 1613
rect 3518 1609 3519 1613
rect 3831 1632 3832 1636
rect 3834 1632 3835 1636
rect 3535 1609 3536 1613
rect 3538 1609 3539 1613
rect 3691 1609 3692 1613
rect 3694 1609 3695 1613
rect 3707 1609 3708 1613
rect 3710 1609 3718 1613
rect 3720 1609 3722 1613
rect 3726 1609 3728 1613
rect 3730 1609 3738 1613
rect 3740 1609 3741 1613
rect 3757 1609 3758 1613
rect 3760 1609 3761 1613
rect 4257 1590 4258 1594
rect 4260 1590 4262 1594
rect 4266 1590 4268 1594
rect 4270 1590 4271 1594
rect 1321 1539 1322 1543
rect 1324 1539 1326 1543
rect 1330 1539 1332 1543
rect 1334 1539 1335 1543
rect 1349 1539 1350 1543
rect 1352 1539 1353 1543
rect 1016 1531 1017 1535
rect 1019 1531 1027 1535
rect 1029 1531 1031 1535
rect 1059 1531 1060 1535
rect 1062 1531 1063 1535
rect 1016 1442 1017 1446
rect 1019 1442 1027 1446
rect 1029 1442 1031 1446
rect 1059 1442 1060 1446
rect 1062 1442 1063 1446
rect 1726 1433 1727 1437
rect 1729 1433 1737 1437
rect 1739 1433 1741 1437
rect 1769 1433 1770 1437
rect 1772 1433 1773 1437
rect 1812 1433 1813 1437
rect 1815 1433 1823 1437
rect 1825 1433 1827 1437
rect 1855 1433 1856 1437
rect 1858 1433 1859 1437
rect 1902 1433 1903 1437
rect 1905 1433 1913 1437
rect 1915 1433 1917 1437
rect 1945 1433 1946 1437
rect 1948 1433 1949 1437
rect 1997 1433 1998 1437
rect 2000 1433 2008 1437
rect 2010 1433 2012 1437
rect 2040 1433 2041 1437
rect 2043 1433 2044 1437
rect 2081 1433 2082 1437
rect 2084 1433 2092 1437
rect 2094 1433 2096 1437
rect 2124 1433 2125 1437
rect 2127 1433 2128 1437
rect 2167 1433 2168 1437
rect 2170 1433 2178 1437
rect 2180 1433 2182 1437
rect 2210 1433 2211 1437
rect 2213 1433 2214 1437
rect 2257 1433 2258 1437
rect 2260 1433 2268 1437
rect 2270 1433 2272 1437
rect 2300 1433 2301 1437
rect 2303 1433 2304 1437
rect 2352 1433 2353 1437
rect 2355 1433 2363 1437
rect 2365 1433 2367 1437
rect 2395 1433 2396 1437
rect 2398 1433 2399 1437
rect 3028 1425 3029 1429
rect 3031 1425 3039 1429
rect 3041 1425 3043 1429
rect 3071 1425 3072 1429
rect 3074 1425 3075 1429
rect 3230 1427 3231 1431
rect 3233 1427 3241 1431
rect 3243 1427 3251 1431
rect 3253 1427 3255 1431
rect 3283 1427 3284 1431
rect 3286 1427 3287 1431
rect 3485 1428 3486 1432
rect 3488 1428 3496 1432
rect 3498 1428 3506 1432
rect 3508 1428 3516 1432
rect 3518 1428 3520 1432
rect 3546 1428 3547 1432
rect 3549 1428 3550 1432
rect 3746 1431 3747 1435
rect 3749 1431 3757 1435
rect 3759 1431 3767 1435
rect 3769 1431 3777 1435
rect 3779 1431 3787 1435
rect 3789 1431 3791 1435
rect 3819 1431 3820 1435
rect 3822 1431 3823 1435
rect 1016 1359 1017 1363
rect 1019 1359 1027 1363
rect 1029 1359 1031 1363
rect 1059 1359 1060 1363
rect 1062 1359 1063 1363
rect 4007 1358 4008 1362
rect 4010 1358 4012 1362
rect 4016 1358 4018 1362
rect 4020 1358 4021 1362
rect 4025 1358 4027 1362
rect 4029 1358 4031 1362
rect 4035 1358 4037 1362
rect 4039 1358 4041 1362
rect 4055 1358 4056 1362
rect 4058 1358 4059 1362
rect 3088 1274 3089 1278
rect 3091 1274 3092 1278
rect 3144 1274 3145 1278
rect 3147 1274 3148 1278
rect 3341 1274 3342 1278
rect 3344 1274 3345 1278
rect 3604 1274 3605 1278
rect 3607 1274 3608 1278
rect 1770 1116 1771 1120
rect 1773 1116 1781 1120
rect 1783 1116 1785 1120
rect 1813 1116 1814 1120
rect 1816 1116 1817 1120
rect 1856 1116 1857 1120
rect 1859 1116 1867 1120
rect 1869 1116 1871 1120
rect 1899 1116 1900 1120
rect 1902 1116 1903 1120
rect 1946 1116 1947 1120
rect 1949 1116 1957 1120
rect 1959 1116 1961 1120
rect 1989 1116 1990 1120
rect 1992 1116 1993 1120
rect 2041 1116 2042 1120
rect 2044 1116 2052 1120
rect 2054 1116 2056 1120
rect 2084 1116 2085 1120
rect 2087 1116 2088 1120
rect 2125 1116 2126 1120
rect 2128 1116 2136 1120
rect 2138 1116 2140 1120
rect 2168 1116 2169 1120
rect 2171 1116 2172 1120
rect 2211 1116 2212 1120
rect 2214 1116 2222 1120
rect 2224 1116 2226 1120
rect 2254 1116 2255 1120
rect 2257 1116 2258 1120
rect 2301 1116 2302 1120
rect 2304 1116 2312 1120
rect 2314 1116 2316 1120
rect 2344 1116 2345 1120
rect 2347 1116 2348 1120
rect 2396 1116 2397 1120
rect 2399 1116 2407 1120
rect 2409 1116 2411 1120
rect 2439 1116 2440 1120
rect 2442 1116 2443 1120
rect 1832 1015 1833 1019
rect 1835 1015 1843 1019
rect 1845 1015 1847 1019
rect 1875 1015 1876 1019
rect 1878 1015 1879 1019
rect 1918 1015 1919 1019
rect 1921 1015 1929 1019
rect 1931 1015 1933 1019
rect 1961 1015 1962 1019
rect 1964 1015 1965 1019
rect 2008 1015 2009 1019
rect 2011 1015 2019 1019
rect 2021 1015 2023 1019
rect 2051 1015 2052 1019
rect 2054 1015 2055 1019
rect 2103 1015 2104 1019
rect 2106 1015 2114 1019
rect 2116 1015 2118 1019
rect 2146 1015 2147 1019
rect 2149 1015 2150 1019
<< pdiffusion >>
rect 1615 3396 1616 3402
rect 1618 3396 1619 3402
rect 1631 3396 1632 3402
rect 1634 3396 1642 3402
rect 1644 3396 1646 3402
rect 1650 3396 1652 3402
rect 1654 3396 1662 3402
rect 1664 3396 1665 3402
rect 1681 3396 1682 3402
rect 1684 3396 1685 3402
rect 1777 3405 1778 3411
rect 1780 3405 1781 3411
rect 1793 3405 1794 3411
rect 1796 3405 1804 3411
rect 1806 3405 1808 3411
rect 1812 3405 1814 3411
rect 1816 3405 1824 3411
rect 1826 3405 1827 3411
rect 1843 3405 1844 3411
rect 1846 3405 1847 3411
rect 2014 3415 2015 3421
rect 2017 3415 2018 3421
rect 2030 3415 2031 3421
rect 2033 3415 2041 3421
rect 2043 3415 2045 3421
rect 2049 3415 2051 3421
rect 2053 3415 2061 3421
rect 2063 3415 2064 3421
rect 2080 3415 2081 3421
rect 2083 3415 2084 3421
rect 1903 3289 1904 3295
rect 1906 3289 1908 3295
rect 1912 3289 1914 3295
rect 1916 3289 1918 3295
rect 1946 3289 1947 3295
rect 1949 3289 1950 3295
rect 2031 3290 2032 3296
rect 2034 3290 2036 3296
rect 2040 3290 2042 3296
rect 2044 3290 2046 3296
rect 2074 3290 2075 3296
rect 2077 3290 2078 3296
rect 2072 3218 2073 3224
rect 2075 3218 2083 3224
rect 2085 3218 2086 3224
rect 2100 3218 2101 3224
rect 2103 3218 2104 3224
rect 1624 3064 1625 3070
rect 1627 3064 1628 3070
rect 1640 3064 1641 3070
rect 1643 3064 1651 3070
rect 1653 3064 1655 3070
rect 1659 3064 1661 3070
rect 1663 3064 1671 3070
rect 1673 3064 1674 3070
rect 1690 3064 1691 3070
rect 1693 3064 1694 3070
rect 1786 3073 1787 3079
rect 1789 3073 1790 3079
rect 1802 3073 1803 3079
rect 1805 3073 1813 3079
rect 1815 3073 1817 3079
rect 1821 3073 1823 3079
rect 1825 3073 1833 3079
rect 1835 3073 1836 3079
rect 1852 3073 1853 3079
rect 1855 3073 1856 3079
rect 2023 3083 2024 3089
rect 2026 3083 2027 3089
rect 2039 3083 2040 3089
rect 2042 3083 2050 3089
rect 2052 3083 2054 3089
rect 2058 3083 2060 3089
rect 2062 3083 2070 3089
rect 2072 3083 2073 3089
rect 2089 3083 2090 3089
rect 2092 3083 2093 3089
rect 1912 2957 1913 2963
rect 1915 2957 1917 2963
rect 1921 2957 1923 2963
rect 1925 2957 1927 2963
rect 1955 2957 1956 2963
rect 1958 2957 1959 2963
rect 2040 2958 2041 2964
rect 2043 2958 2045 2964
rect 2049 2958 2051 2964
rect 2053 2958 2055 2964
rect 2083 2958 2084 2964
rect 2086 2958 2087 2964
rect 2081 2886 2082 2892
rect 2084 2886 2092 2892
rect 2094 2886 2095 2892
rect 2109 2886 2110 2892
rect 2112 2886 2113 2892
rect 1645 2698 1646 2704
rect 1648 2698 1649 2704
rect 1661 2698 1662 2704
rect 1664 2698 1672 2704
rect 1674 2698 1676 2704
rect 1680 2698 1682 2704
rect 1684 2698 1692 2704
rect 1694 2698 1695 2704
rect 1711 2698 1712 2704
rect 1714 2698 1715 2704
rect 1807 2707 1808 2713
rect 1810 2707 1811 2713
rect 1823 2707 1824 2713
rect 1826 2707 1834 2713
rect 1836 2707 1838 2713
rect 1842 2707 1844 2713
rect 1846 2707 1854 2713
rect 1856 2707 1857 2713
rect 1873 2707 1874 2713
rect 1876 2707 1877 2713
rect 2044 2717 2045 2723
rect 2047 2717 2048 2723
rect 2060 2717 2061 2723
rect 2063 2717 2071 2723
rect 2073 2717 2075 2723
rect 2079 2717 2081 2723
rect 2083 2717 2091 2723
rect 2093 2717 2094 2723
rect 2110 2717 2111 2723
rect 2113 2717 2114 2723
rect 1933 2591 1934 2597
rect 1936 2591 1938 2597
rect 1942 2591 1944 2597
rect 1946 2591 1948 2597
rect 1976 2591 1977 2597
rect 1979 2591 1980 2597
rect 2061 2592 2062 2598
rect 2064 2592 2066 2598
rect 2070 2592 2072 2598
rect 2074 2592 2076 2598
rect 2104 2592 2105 2598
rect 2107 2592 2108 2598
rect 2102 2520 2103 2526
rect 2105 2520 2113 2526
rect 2115 2520 2116 2526
rect 2130 2520 2131 2526
rect 2133 2520 2134 2526
rect 1673 2324 1674 2330
rect 1676 2324 1677 2330
rect 1689 2324 1690 2330
rect 1692 2324 1700 2330
rect 1702 2324 1704 2330
rect 1708 2324 1710 2330
rect 1712 2324 1720 2330
rect 1722 2324 1723 2330
rect 1739 2324 1740 2330
rect 1742 2324 1743 2330
rect 1835 2333 1836 2339
rect 1838 2333 1839 2339
rect 1851 2333 1852 2339
rect 1854 2333 1862 2339
rect 1864 2333 1866 2339
rect 1870 2333 1872 2339
rect 1874 2333 1882 2339
rect 1884 2333 1885 2339
rect 1901 2333 1902 2339
rect 1904 2333 1905 2339
rect 2072 2343 2073 2349
rect 2075 2343 2076 2349
rect 2088 2343 2089 2349
rect 2091 2343 2099 2349
rect 2101 2343 2103 2349
rect 2107 2343 2109 2349
rect 2111 2343 2119 2349
rect 2121 2343 2122 2349
rect 2138 2343 2139 2349
rect 2141 2343 2142 2349
rect 1961 2217 1962 2223
rect 1964 2217 1966 2223
rect 1970 2217 1972 2223
rect 1974 2217 1976 2223
rect 2004 2217 2005 2223
rect 2007 2217 2008 2223
rect 2089 2218 2090 2224
rect 2092 2218 2094 2224
rect 2098 2218 2100 2224
rect 2102 2218 2104 2224
rect 2132 2218 2133 2224
rect 2135 2218 2136 2224
rect 2130 2146 2131 2152
rect 2133 2146 2141 2152
rect 2143 2146 2144 2152
rect 2158 2146 2159 2152
rect 2161 2146 2162 2152
rect 3958 1781 3959 1787
rect 3961 1781 3963 1787
rect 3967 1781 3969 1787
rect 3971 1781 3973 1787
rect 3977 1781 3979 1787
rect 3981 1781 3983 1787
rect 3987 1781 3989 1787
rect 3991 1781 3993 1787
rect 4019 1781 4020 1787
rect 4022 1781 4023 1787
rect 1052 1723 1053 1727
rect 1055 1723 1056 1727
rect 1108 1723 1109 1727
rect 1111 1723 1112 1727
rect 1748 1707 1749 1713
rect 1751 1707 1753 1713
rect 1757 1707 1759 1713
rect 1761 1707 1763 1713
rect 1791 1707 1792 1713
rect 1794 1707 1795 1713
rect 1834 1707 1835 1713
rect 1837 1707 1839 1713
rect 1843 1707 1845 1713
rect 1847 1707 1849 1713
rect 1877 1707 1878 1713
rect 1880 1707 1881 1713
rect 1924 1707 1925 1713
rect 1927 1707 1929 1713
rect 1933 1707 1935 1713
rect 1937 1707 1939 1713
rect 1967 1707 1968 1713
rect 1970 1707 1971 1713
rect 2019 1707 2020 1713
rect 2022 1707 2024 1713
rect 2028 1707 2030 1713
rect 2032 1707 2034 1713
rect 2062 1707 2063 1713
rect 2065 1707 2066 1713
rect 2103 1707 2104 1713
rect 2106 1707 2108 1713
rect 2112 1707 2114 1713
rect 2116 1707 2118 1713
rect 2146 1707 2147 1713
rect 2149 1707 2150 1713
rect 2189 1707 2190 1713
rect 2192 1707 2194 1713
rect 2198 1707 2200 1713
rect 2202 1707 2204 1713
rect 2232 1707 2233 1713
rect 2235 1707 2236 1713
rect 2279 1707 2280 1713
rect 2282 1707 2284 1713
rect 2288 1707 2290 1713
rect 2292 1707 2294 1713
rect 2322 1707 2323 1713
rect 2325 1707 2326 1713
rect 2374 1707 2375 1713
rect 2377 1707 2379 1713
rect 2383 1707 2385 1713
rect 2387 1707 2389 1713
rect 2417 1707 2418 1713
rect 2420 1707 2421 1713
rect 2963 1655 2964 1661
rect 2966 1655 2967 1661
rect 2979 1655 2980 1661
rect 2982 1655 2990 1661
rect 2992 1655 2994 1661
rect 2998 1655 3000 1661
rect 3002 1655 3010 1661
rect 3012 1655 3013 1661
rect 3029 1655 3030 1661
rect 3032 1655 3033 1661
rect 1015 1646 1016 1652
rect 1018 1646 1020 1652
rect 1024 1646 1026 1652
rect 1028 1646 1030 1652
rect 1058 1646 1059 1652
rect 1061 1646 1062 1652
rect 3103 1652 3104 1656
rect 3106 1652 3107 1656
rect 3212 1655 3213 1661
rect 3215 1655 3216 1661
rect 3228 1655 3229 1661
rect 3231 1655 3239 1661
rect 3241 1655 3243 1661
rect 3247 1655 3249 1661
rect 3251 1655 3259 1661
rect 3261 1655 3262 1661
rect 3278 1655 3279 1661
rect 3281 1655 3282 1661
rect 3352 1652 3353 1656
rect 3355 1652 3356 1656
rect 3469 1655 3470 1661
rect 3472 1655 3473 1661
rect 3485 1655 3486 1661
rect 3488 1655 3496 1661
rect 3498 1655 3500 1661
rect 3504 1655 3506 1661
rect 3508 1655 3516 1661
rect 3518 1655 3519 1661
rect 3535 1655 3536 1661
rect 3538 1655 3539 1661
rect 3609 1652 3610 1656
rect 3612 1652 3613 1656
rect 3691 1655 3692 1661
rect 3694 1655 3695 1661
rect 3707 1655 3708 1661
rect 3710 1655 3718 1661
rect 3720 1655 3722 1661
rect 3726 1655 3728 1661
rect 3730 1655 3738 1661
rect 3740 1655 3741 1661
rect 3757 1655 3758 1661
rect 3760 1655 3761 1661
rect 3831 1652 3832 1656
rect 3834 1652 3835 1656
rect 4257 1626 4258 1632
rect 4260 1626 4268 1632
rect 4270 1626 4271 1632
rect 1321 1575 1322 1581
rect 1324 1575 1332 1581
rect 1334 1575 1335 1581
rect 1349 1575 1350 1581
rect 1352 1575 1353 1581
rect 1016 1561 1017 1567
rect 1019 1561 1021 1567
rect 1025 1561 1027 1567
rect 1029 1561 1031 1567
rect 1059 1561 1060 1567
rect 1062 1561 1063 1567
rect 1016 1472 1017 1478
rect 1019 1472 1021 1478
rect 1025 1472 1027 1478
rect 1029 1472 1031 1478
rect 1059 1472 1060 1478
rect 1062 1472 1063 1478
rect 3746 1479 3747 1485
rect 3749 1479 3751 1485
rect 3755 1479 3757 1485
rect 3759 1479 3761 1485
rect 3765 1479 3767 1485
rect 3769 1479 3771 1485
rect 3775 1479 3777 1485
rect 3779 1479 3781 1485
rect 3785 1479 3787 1485
rect 3789 1479 3791 1485
rect 3819 1479 3820 1485
rect 3822 1479 3823 1485
rect 1726 1463 1727 1469
rect 1729 1463 1731 1469
rect 1735 1463 1737 1469
rect 1739 1463 1741 1469
rect 1769 1463 1770 1469
rect 1772 1463 1773 1469
rect 1812 1463 1813 1469
rect 1815 1463 1817 1469
rect 1821 1463 1823 1469
rect 1825 1463 1827 1469
rect 1855 1463 1856 1469
rect 1858 1463 1859 1469
rect 1902 1463 1903 1469
rect 1905 1463 1907 1469
rect 1911 1463 1913 1469
rect 1915 1463 1917 1469
rect 1945 1463 1946 1469
rect 1948 1463 1949 1469
rect 1997 1463 1998 1469
rect 2000 1463 2002 1469
rect 2006 1463 2008 1469
rect 2010 1463 2012 1469
rect 2040 1463 2041 1469
rect 2043 1463 2044 1469
rect 2081 1463 2082 1469
rect 2084 1463 2086 1469
rect 2090 1463 2092 1469
rect 2094 1463 2096 1469
rect 2124 1463 2125 1469
rect 2127 1463 2128 1469
rect 2167 1463 2168 1469
rect 2170 1463 2172 1469
rect 2176 1463 2178 1469
rect 2180 1463 2182 1469
rect 2210 1463 2211 1469
rect 2213 1463 2214 1469
rect 2257 1463 2258 1469
rect 2260 1463 2262 1469
rect 2266 1463 2268 1469
rect 2270 1463 2272 1469
rect 2300 1463 2301 1469
rect 2303 1463 2304 1469
rect 2352 1463 2353 1469
rect 2355 1463 2357 1469
rect 2361 1463 2363 1469
rect 2365 1463 2367 1469
rect 2395 1463 2396 1469
rect 2398 1463 2399 1469
rect 3485 1469 3486 1475
rect 3488 1469 3490 1475
rect 3494 1469 3496 1475
rect 3498 1469 3500 1475
rect 3504 1469 3506 1475
rect 3508 1469 3510 1475
rect 3514 1469 3516 1475
rect 3518 1469 3520 1475
rect 3546 1469 3547 1475
rect 3549 1469 3550 1475
rect 3028 1455 3029 1461
rect 3031 1455 3033 1461
rect 3037 1455 3039 1461
rect 3041 1455 3043 1461
rect 3071 1455 3072 1461
rect 3074 1455 3075 1461
rect 3230 1460 3231 1466
rect 3233 1460 3235 1466
rect 3239 1460 3241 1466
rect 3243 1460 3245 1466
rect 3249 1460 3251 1466
rect 3253 1460 3255 1466
rect 3283 1460 3284 1466
rect 3286 1460 3287 1466
rect 4007 1408 4008 1414
rect 4010 1408 4018 1414
rect 4020 1408 4027 1414
rect 4029 1408 4037 1414
rect 4039 1408 4041 1414
rect 4055 1408 4056 1414
rect 4058 1408 4059 1414
rect 1016 1389 1017 1395
rect 1019 1389 1021 1395
rect 1025 1389 1027 1395
rect 1029 1389 1031 1395
rect 1059 1389 1060 1395
rect 1062 1389 1063 1395
rect 3088 1294 3089 1298
rect 3091 1294 3092 1298
rect 3144 1294 3145 1298
rect 3147 1294 3148 1298
rect 3341 1294 3342 1298
rect 3344 1294 3345 1298
rect 3604 1294 3605 1298
rect 3607 1294 3608 1298
rect 1770 1146 1771 1152
rect 1773 1146 1775 1152
rect 1779 1146 1781 1152
rect 1783 1146 1785 1152
rect 1813 1146 1814 1152
rect 1816 1146 1817 1152
rect 1856 1146 1857 1152
rect 1859 1146 1861 1152
rect 1865 1146 1867 1152
rect 1869 1146 1871 1152
rect 1899 1146 1900 1152
rect 1902 1146 1903 1152
rect 1946 1146 1947 1152
rect 1949 1146 1951 1152
rect 1955 1146 1957 1152
rect 1959 1146 1961 1152
rect 1989 1146 1990 1152
rect 1992 1146 1993 1152
rect 2041 1146 2042 1152
rect 2044 1146 2046 1152
rect 2050 1146 2052 1152
rect 2054 1146 2056 1152
rect 2084 1146 2085 1152
rect 2087 1146 2088 1152
rect 2125 1146 2126 1152
rect 2128 1146 2130 1152
rect 2134 1146 2136 1152
rect 2138 1146 2140 1152
rect 2168 1146 2169 1152
rect 2171 1146 2172 1152
rect 2211 1146 2212 1152
rect 2214 1146 2216 1152
rect 2220 1146 2222 1152
rect 2224 1146 2226 1152
rect 2254 1146 2255 1152
rect 2257 1146 2258 1152
rect 2301 1146 2302 1152
rect 2304 1146 2306 1152
rect 2310 1146 2312 1152
rect 2314 1146 2316 1152
rect 2344 1146 2345 1152
rect 2347 1146 2348 1152
rect 2396 1146 2397 1152
rect 2399 1146 2401 1152
rect 2405 1146 2407 1152
rect 2409 1146 2411 1152
rect 2439 1146 2440 1152
rect 2442 1146 2443 1152
rect 1832 1045 1833 1051
rect 1835 1045 1837 1051
rect 1841 1045 1843 1051
rect 1845 1045 1847 1051
rect 1875 1045 1876 1051
rect 1878 1045 1879 1051
rect 1918 1045 1919 1051
rect 1921 1045 1923 1051
rect 1927 1045 1929 1051
rect 1931 1045 1933 1051
rect 1961 1045 1962 1051
rect 1964 1045 1965 1051
rect 2008 1045 2009 1051
rect 2011 1045 2013 1051
rect 2017 1045 2019 1051
rect 2021 1045 2023 1051
rect 2051 1045 2052 1051
rect 2054 1045 2055 1051
rect 2103 1045 2104 1051
rect 2106 1045 2108 1051
rect 2112 1045 2114 1051
rect 2116 1045 2118 1051
rect 2146 1045 2147 1051
rect 2149 1045 2150 1051
<< ndcontact >>
rect 1611 3350 1615 3354
rect 1619 3350 1623 3354
rect 1627 3350 1631 3354
rect 1646 3350 1650 3354
rect 1665 3350 1669 3354
rect 1773 3359 1777 3363
rect 1781 3359 1785 3363
rect 1789 3359 1793 3363
rect 1808 3359 1812 3363
rect 1827 3359 1831 3363
rect 1677 3350 1681 3354
rect 1685 3350 1689 3354
rect 2010 3369 2014 3373
rect 2018 3369 2022 3373
rect 2026 3369 2030 3373
rect 2045 3369 2049 3373
rect 2064 3369 2068 3373
rect 1839 3359 1843 3363
rect 1847 3359 1851 3363
rect 2076 3369 2080 3373
rect 2084 3369 2088 3373
rect 1899 3259 1903 3263
rect 1918 3259 1922 3263
rect 1942 3259 1946 3263
rect 1950 3259 1954 3263
rect 2027 3260 2031 3264
rect 2046 3260 2050 3264
rect 2070 3260 2074 3264
rect 2078 3260 2082 3264
rect 2068 3182 2072 3186
rect 2077 3182 2081 3186
rect 2086 3182 2090 3186
rect 2096 3182 2100 3186
rect 2104 3182 2108 3186
rect 1620 3018 1624 3022
rect 1628 3018 1632 3022
rect 1636 3018 1640 3022
rect 1655 3018 1659 3022
rect 1674 3018 1678 3022
rect 1782 3027 1786 3031
rect 1790 3027 1794 3031
rect 1798 3027 1802 3031
rect 1817 3027 1821 3031
rect 1836 3027 1840 3031
rect 1686 3018 1690 3022
rect 1694 3018 1698 3022
rect 2019 3037 2023 3041
rect 2027 3037 2031 3041
rect 2035 3037 2039 3041
rect 2054 3037 2058 3041
rect 2073 3037 2077 3041
rect 1848 3027 1852 3031
rect 1856 3027 1860 3031
rect 2085 3037 2089 3041
rect 2093 3037 2097 3041
rect 1908 2927 1912 2931
rect 1927 2927 1931 2931
rect 1951 2927 1955 2931
rect 1959 2927 1963 2931
rect 2036 2928 2040 2932
rect 2055 2928 2059 2932
rect 2079 2928 2083 2932
rect 2087 2928 2091 2932
rect 2077 2850 2081 2854
rect 2086 2850 2090 2854
rect 2095 2850 2099 2854
rect 2105 2850 2109 2854
rect 2113 2850 2117 2854
rect 1641 2652 1645 2656
rect 1649 2652 1653 2656
rect 1657 2652 1661 2656
rect 1676 2652 1680 2656
rect 1695 2652 1699 2656
rect 1803 2661 1807 2665
rect 1811 2661 1815 2665
rect 1819 2661 1823 2665
rect 1838 2661 1842 2665
rect 1857 2661 1861 2665
rect 1707 2652 1711 2656
rect 1715 2652 1719 2656
rect 2040 2671 2044 2675
rect 2048 2671 2052 2675
rect 2056 2671 2060 2675
rect 2075 2671 2079 2675
rect 2094 2671 2098 2675
rect 1869 2661 1873 2665
rect 1877 2661 1881 2665
rect 2106 2671 2110 2675
rect 2114 2671 2118 2675
rect 1929 2561 1933 2565
rect 1948 2561 1952 2565
rect 1972 2561 1976 2565
rect 1980 2561 1984 2565
rect 2057 2562 2061 2566
rect 2076 2562 2080 2566
rect 2100 2562 2104 2566
rect 2108 2562 2112 2566
rect 2098 2484 2102 2488
rect 2107 2484 2111 2488
rect 2116 2484 2120 2488
rect 2126 2484 2130 2488
rect 2134 2484 2138 2488
rect 1669 2278 1673 2282
rect 1677 2278 1681 2282
rect 1685 2278 1689 2282
rect 1704 2278 1708 2282
rect 1723 2278 1727 2282
rect 1831 2287 1835 2291
rect 1839 2287 1843 2291
rect 1847 2287 1851 2291
rect 1866 2287 1870 2291
rect 1885 2287 1889 2291
rect 1735 2278 1739 2282
rect 1743 2278 1747 2282
rect 2068 2297 2072 2301
rect 2076 2297 2080 2301
rect 2084 2297 2088 2301
rect 2103 2297 2107 2301
rect 2122 2297 2126 2301
rect 1897 2287 1901 2291
rect 1905 2287 1909 2291
rect 2134 2297 2138 2301
rect 2142 2297 2146 2301
rect 1957 2187 1961 2191
rect 1976 2187 1980 2191
rect 2000 2187 2004 2191
rect 2008 2187 2012 2191
rect 2085 2188 2089 2192
rect 2104 2188 2108 2192
rect 2128 2188 2132 2192
rect 2136 2188 2140 2192
rect 2126 2110 2130 2114
rect 2135 2110 2139 2114
rect 2144 2110 2148 2114
rect 2154 2110 2158 2114
rect 2162 2110 2166 2114
rect 3954 1740 3958 1744
rect 3993 1740 3997 1744
rect 4015 1740 4019 1744
rect 4023 1740 4027 1744
rect 1048 1703 1052 1707
rect 1056 1703 1060 1707
rect 1104 1703 1108 1707
rect 1112 1703 1116 1707
rect 1744 1677 1748 1681
rect 1763 1677 1767 1681
rect 1787 1677 1791 1681
rect 1795 1677 1799 1681
rect 1830 1677 1834 1681
rect 1849 1677 1853 1681
rect 1873 1677 1877 1681
rect 1881 1677 1885 1681
rect 1920 1677 1924 1681
rect 1939 1677 1943 1681
rect 1963 1677 1967 1681
rect 1971 1677 1975 1681
rect 2015 1677 2019 1681
rect 2034 1677 2038 1681
rect 2058 1677 2062 1681
rect 2066 1677 2070 1681
rect 2099 1677 2103 1681
rect 2118 1677 2122 1681
rect 2142 1677 2146 1681
rect 2150 1677 2154 1681
rect 2185 1677 2189 1681
rect 2204 1677 2208 1681
rect 2228 1677 2232 1681
rect 2236 1677 2240 1681
rect 2275 1677 2279 1681
rect 2294 1677 2298 1681
rect 2318 1677 2322 1681
rect 2326 1677 2330 1681
rect 2370 1677 2374 1681
rect 2389 1677 2393 1681
rect 2413 1677 2417 1681
rect 2421 1677 2425 1681
rect 1011 1616 1015 1620
rect 1030 1616 1034 1620
rect 1054 1616 1058 1620
rect 1062 1616 1066 1620
rect 3099 1632 3103 1636
rect 3107 1632 3111 1636
rect 2959 1609 2963 1613
rect 2967 1609 2971 1613
rect 2975 1609 2979 1613
rect 2994 1609 2998 1613
rect 3013 1609 3017 1613
rect 3348 1632 3352 1636
rect 3356 1632 3360 1636
rect 3025 1609 3029 1613
rect 3033 1609 3037 1613
rect 3208 1609 3212 1613
rect 3216 1609 3220 1613
rect 3224 1609 3228 1613
rect 3243 1609 3247 1613
rect 3262 1609 3266 1613
rect 3605 1632 3609 1636
rect 3613 1632 3617 1636
rect 3274 1609 3278 1613
rect 3282 1609 3286 1613
rect 3465 1609 3469 1613
rect 3473 1609 3477 1613
rect 3481 1609 3485 1613
rect 3500 1609 3504 1613
rect 3519 1609 3523 1613
rect 3827 1632 3831 1636
rect 3835 1632 3839 1636
rect 3531 1609 3535 1613
rect 3539 1609 3543 1613
rect 3687 1609 3691 1613
rect 3695 1609 3699 1613
rect 3703 1609 3707 1613
rect 3722 1609 3726 1613
rect 3741 1609 3745 1613
rect 3753 1609 3757 1613
rect 3761 1609 3765 1613
rect 4253 1590 4257 1594
rect 4262 1590 4266 1594
rect 4271 1590 4275 1594
rect 1317 1539 1321 1543
rect 1326 1539 1330 1543
rect 1335 1539 1339 1543
rect 1345 1539 1349 1543
rect 1353 1539 1357 1543
rect 1012 1531 1016 1535
rect 1031 1531 1035 1535
rect 1055 1531 1059 1535
rect 1063 1531 1067 1535
rect 1012 1442 1016 1446
rect 1031 1442 1035 1446
rect 1055 1442 1059 1446
rect 1063 1442 1067 1446
rect 1722 1433 1726 1437
rect 1741 1433 1745 1437
rect 1765 1433 1769 1437
rect 1773 1433 1777 1437
rect 1808 1433 1812 1437
rect 1827 1433 1831 1437
rect 1851 1433 1855 1437
rect 1859 1433 1863 1437
rect 1898 1433 1902 1437
rect 1917 1433 1921 1437
rect 1941 1433 1945 1437
rect 1949 1433 1953 1437
rect 1993 1433 1997 1437
rect 2012 1433 2016 1437
rect 2036 1433 2040 1437
rect 2044 1433 2048 1437
rect 2077 1433 2081 1437
rect 2096 1433 2100 1437
rect 2120 1433 2124 1437
rect 2128 1433 2132 1437
rect 2163 1433 2167 1437
rect 2182 1433 2186 1437
rect 2206 1433 2210 1437
rect 2214 1433 2218 1437
rect 2253 1433 2257 1437
rect 2272 1433 2276 1437
rect 2296 1433 2300 1437
rect 2304 1433 2308 1437
rect 2348 1433 2352 1437
rect 2367 1433 2371 1437
rect 2391 1433 2395 1437
rect 2399 1433 2403 1437
rect 3024 1425 3028 1429
rect 3043 1425 3047 1429
rect 3067 1425 3071 1429
rect 3075 1425 3079 1429
rect 3226 1427 3230 1431
rect 3255 1427 3259 1431
rect 3279 1427 3283 1431
rect 3287 1427 3291 1431
rect 3481 1428 3485 1432
rect 3520 1428 3524 1432
rect 3542 1428 3546 1432
rect 3550 1428 3554 1432
rect 3742 1431 3746 1435
rect 3791 1431 3795 1435
rect 3815 1431 3819 1435
rect 3823 1431 3827 1435
rect 1012 1359 1016 1363
rect 1031 1359 1035 1363
rect 1055 1359 1059 1363
rect 1063 1359 1067 1363
rect 4003 1358 4007 1362
rect 4012 1358 4016 1362
rect 4021 1358 4025 1362
rect 4031 1358 4035 1362
rect 4041 1358 4045 1362
rect 4051 1358 4055 1362
rect 4059 1358 4063 1362
rect 3084 1274 3088 1278
rect 3092 1274 3096 1278
rect 3140 1274 3144 1278
rect 3148 1274 3152 1278
rect 3337 1274 3341 1278
rect 3345 1274 3349 1278
rect 3600 1274 3604 1278
rect 3608 1274 3612 1278
rect 1766 1116 1770 1120
rect 1785 1116 1789 1120
rect 1809 1116 1813 1120
rect 1817 1116 1821 1120
rect 1852 1116 1856 1120
rect 1871 1116 1875 1120
rect 1895 1116 1899 1120
rect 1903 1116 1907 1120
rect 1942 1116 1946 1120
rect 1961 1116 1965 1120
rect 1985 1116 1989 1120
rect 1993 1116 1997 1120
rect 2037 1116 2041 1120
rect 2056 1116 2060 1120
rect 2080 1116 2084 1120
rect 2088 1116 2092 1120
rect 2121 1116 2125 1120
rect 2140 1116 2144 1120
rect 2164 1116 2168 1120
rect 2172 1116 2176 1120
rect 2207 1116 2211 1120
rect 2226 1116 2230 1120
rect 2250 1116 2254 1120
rect 2258 1116 2262 1120
rect 2297 1116 2301 1120
rect 2316 1116 2320 1120
rect 2340 1116 2344 1120
rect 2348 1116 2352 1120
rect 2392 1116 2396 1120
rect 2411 1116 2415 1120
rect 2435 1116 2439 1120
rect 2443 1116 2447 1120
rect 1828 1015 1832 1019
rect 1847 1015 1851 1019
rect 1871 1015 1875 1019
rect 1879 1015 1883 1019
rect 1914 1015 1918 1019
rect 1933 1015 1937 1019
rect 1957 1015 1961 1019
rect 1965 1015 1969 1019
rect 2004 1015 2008 1019
rect 2023 1015 2027 1019
rect 2047 1015 2051 1019
rect 2055 1015 2059 1019
rect 2099 1015 2103 1019
rect 2118 1015 2122 1019
rect 2142 1015 2146 1019
rect 2150 1015 2154 1019
<< pdcontact >>
rect 1611 3396 1615 3402
rect 1619 3396 1623 3402
rect 1627 3396 1631 3402
rect 1646 3396 1650 3402
rect 1665 3396 1669 3402
rect 1677 3396 1681 3402
rect 1685 3396 1689 3402
rect 1773 3405 1777 3411
rect 1781 3405 1785 3411
rect 1789 3405 1793 3411
rect 1808 3405 1812 3411
rect 1827 3405 1831 3411
rect 1839 3405 1843 3411
rect 1847 3405 1851 3411
rect 2010 3415 2014 3421
rect 2018 3415 2022 3421
rect 2026 3415 2030 3421
rect 2045 3415 2049 3421
rect 2064 3415 2068 3421
rect 2076 3415 2080 3421
rect 2084 3415 2088 3421
rect 1899 3289 1903 3295
rect 1908 3289 1912 3295
rect 1918 3289 1922 3295
rect 1942 3289 1946 3295
rect 1950 3289 1954 3295
rect 2027 3290 2031 3296
rect 2036 3290 2040 3296
rect 2046 3290 2050 3296
rect 2070 3290 2074 3296
rect 2078 3290 2082 3296
rect 2068 3218 2072 3224
rect 2086 3218 2090 3224
rect 2096 3218 2100 3224
rect 2104 3218 2108 3224
rect 1620 3064 1624 3070
rect 1628 3064 1632 3070
rect 1636 3064 1640 3070
rect 1655 3064 1659 3070
rect 1674 3064 1678 3070
rect 1686 3064 1690 3070
rect 1694 3064 1698 3070
rect 1782 3073 1786 3079
rect 1790 3073 1794 3079
rect 1798 3073 1802 3079
rect 1817 3073 1821 3079
rect 1836 3073 1840 3079
rect 1848 3073 1852 3079
rect 1856 3073 1860 3079
rect 2019 3083 2023 3089
rect 2027 3083 2031 3089
rect 2035 3083 2039 3089
rect 2054 3083 2058 3089
rect 2073 3083 2077 3089
rect 2085 3083 2089 3089
rect 2093 3083 2097 3089
rect 1908 2957 1912 2963
rect 1917 2957 1921 2963
rect 1927 2957 1931 2963
rect 1951 2957 1955 2963
rect 1959 2957 1963 2963
rect 2036 2958 2040 2964
rect 2045 2958 2049 2964
rect 2055 2958 2059 2964
rect 2079 2958 2083 2964
rect 2087 2958 2091 2964
rect 2077 2886 2081 2892
rect 2095 2886 2099 2892
rect 2105 2886 2109 2892
rect 2113 2886 2117 2892
rect 1641 2698 1645 2704
rect 1649 2698 1653 2704
rect 1657 2698 1661 2704
rect 1676 2698 1680 2704
rect 1695 2698 1699 2704
rect 1707 2698 1711 2704
rect 1715 2698 1719 2704
rect 1803 2707 1807 2713
rect 1811 2707 1815 2713
rect 1819 2707 1823 2713
rect 1838 2707 1842 2713
rect 1857 2707 1861 2713
rect 1869 2707 1873 2713
rect 1877 2707 1881 2713
rect 2040 2717 2044 2723
rect 2048 2717 2052 2723
rect 2056 2717 2060 2723
rect 2075 2717 2079 2723
rect 2094 2717 2098 2723
rect 2106 2717 2110 2723
rect 2114 2717 2118 2723
rect 1929 2591 1933 2597
rect 1938 2591 1942 2597
rect 1948 2591 1952 2597
rect 1972 2591 1976 2597
rect 1980 2591 1984 2597
rect 2057 2592 2061 2598
rect 2066 2592 2070 2598
rect 2076 2592 2080 2598
rect 2100 2592 2104 2598
rect 2108 2592 2112 2598
rect 2098 2520 2102 2526
rect 2116 2520 2120 2526
rect 2126 2520 2130 2526
rect 2134 2520 2138 2526
rect 1669 2324 1673 2330
rect 1677 2324 1681 2330
rect 1685 2324 1689 2330
rect 1704 2324 1708 2330
rect 1723 2324 1727 2330
rect 1735 2324 1739 2330
rect 1743 2324 1747 2330
rect 1831 2333 1835 2339
rect 1839 2333 1843 2339
rect 1847 2333 1851 2339
rect 1866 2333 1870 2339
rect 1885 2333 1889 2339
rect 1897 2333 1901 2339
rect 1905 2333 1909 2339
rect 2068 2343 2072 2349
rect 2076 2343 2080 2349
rect 2084 2343 2088 2349
rect 2103 2343 2107 2349
rect 2122 2343 2126 2349
rect 2134 2343 2138 2349
rect 2142 2343 2146 2349
rect 1957 2217 1961 2223
rect 1966 2217 1970 2223
rect 1976 2217 1980 2223
rect 2000 2217 2004 2223
rect 2008 2217 2012 2223
rect 2085 2218 2089 2224
rect 2094 2218 2098 2224
rect 2104 2218 2108 2224
rect 2128 2218 2132 2224
rect 2136 2218 2140 2224
rect 2126 2146 2130 2152
rect 2144 2146 2148 2152
rect 2154 2146 2158 2152
rect 2162 2146 2166 2152
rect 3954 1781 3958 1787
rect 3963 1781 3967 1787
rect 3973 1781 3977 1787
rect 3983 1781 3987 1787
rect 3993 1781 3997 1787
rect 4015 1781 4019 1787
rect 4023 1781 4027 1787
rect 1048 1723 1052 1727
rect 1056 1723 1060 1727
rect 1104 1723 1108 1727
rect 1112 1723 1116 1727
rect 1744 1707 1748 1713
rect 1753 1707 1757 1713
rect 1763 1707 1767 1713
rect 1787 1707 1791 1713
rect 1795 1707 1799 1713
rect 1830 1707 1834 1713
rect 1839 1707 1843 1713
rect 1849 1707 1853 1713
rect 1873 1707 1877 1713
rect 1881 1707 1885 1713
rect 1920 1707 1924 1713
rect 1929 1707 1933 1713
rect 1939 1707 1943 1713
rect 1963 1707 1967 1713
rect 1971 1707 1975 1713
rect 2015 1707 2019 1713
rect 2024 1707 2028 1713
rect 2034 1707 2038 1713
rect 2058 1707 2062 1713
rect 2066 1707 2070 1713
rect 2099 1707 2103 1713
rect 2108 1707 2112 1713
rect 2118 1707 2122 1713
rect 2142 1707 2146 1713
rect 2150 1707 2154 1713
rect 2185 1707 2189 1713
rect 2194 1707 2198 1713
rect 2204 1707 2208 1713
rect 2228 1707 2232 1713
rect 2236 1707 2240 1713
rect 2275 1707 2279 1713
rect 2284 1707 2288 1713
rect 2294 1707 2298 1713
rect 2318 1707 2322 1713
rect 2326 1707 2330 1713
rect 2370 1707 2374 1713
rect 2379 1707 2383 1713
rect 2389 1707 2393 1713
rect 2413 1707 2417 1713
rect 2421 1707 2425 1713
rect 2959 1655 2963 1661
rect 2967 1655 2971 1661
rect 2975 1655 2979 1661
rect 2994 1655 2998 1661
rect 3013 1655 3017 1661
rect 3025 1655 3029 1661
rect 3033 1655 3037 1661
rect 1011 1646 1015 1652
rect 1020 1646 1024 1652
rect 1030 1646 1034 1652
rect 1054 1646 1058 1652
rect 1062 1646 1066 1652
rect 3099 1652 3103 1656
rect 3107 1652 3111 1656
rect 3208 1655 3212 1661
rect 3216 1655 3220 1661
rect 3224 1655 3228 1661
rect 3243 1655 3247 1661
rect 3262 1655 3266 1661
rect 3274 1655 3278 1661
rect 3282 1655 3286 1661
rect 3348 1652 3352 1656
rect 3356 1652 3360 1656
rect 3465 1655 3469 1661
rect 3473 1655 3477 1661
rect 3481 1655 3485 1661
rect 3500 1655 3504 1661
rect 3519 1655 3523 1661
rect 3531 1655 3535 1661
rect 3539 1655 3543 1661
rect 3605 1652 3609 1656
rect 3613 1652 3617 1656
rect 3687 1655 3691 1661
rect 3695 1655 3699 1661
rect 3703 1655 3707 1661
rect 3722 1655 3726 1661
rect 3741 1655 3745 1661
rect 3753 1655 3757 1661
rect 3761 1655 3765 1661
rect 3827 1652 3831 1656
rect 3835 1652 3839 1656
rect 4253 1626 4257 1632
rect 4271 1626 4275 1632
rect 1317 1575 1321 1581
rect 1335 1575 1339 1581
rect 1345 1575 1349 1581
rect 1353 1575 1357 1581
rect 1012 1561 1016 1567
rect 1021 1561 1025 1567
rect 1031 1561 1035 1567
rect 1055 1561 1059 1567
rect 1063 1561 1067 1567
rect 1012 1472 1016 1478
rect 1021 1472 1025 1478
rect 1031 1472 1035 1478
rect 1055 1472 1059 1478
rect 1063 1472 1067 1478
rect 3742 1479 3746 1485
rect 3751 1479 3755 1485
rect 3761 1479 3765 1485
rect 3771 1479 3775 1485
rect 3781 1479 3785 1485
rect 3791 1479 3795 1485
rect 3815 1479 3819 1485
rect 3823 1479 3827 1485
rect 1722 1463 1726 1469
rect 1731 1463 1735 1469
rect 1741 1463 1745 1469
rect 1765 1463 1769 1469
rect 1773 1463 1777 1469
rect 1808 1463 1812 1469
rect 1817 1463 1821 1469
rect 1827 1463 1831 1469
rect 1851 1463 1855 1469
rect 1859 1463 1863 1469
rect 1898 1463 1902 1469
rect 1907 1463 1911 1469
rect 1917 1463 1921 1469
rect 1941 1463 1945 1469
rect 1949 1463 1953 1469
rect 1993 1463 1997 1469
rect 2002 1463 2006 1469
rect 2012 1463 2016 1469
rect 2036 1463 2040 1469
rect 2044 1463 2048 1469
rect 2077 1463 2081 1469
rect 2086 1463 2090 1469
rect 2096 1463 2100 1469
rect 2120 1463 2124 1469
rect 2128 1463 2132 1469
rect 2163 1463 2167 1469
rect 2172 1463 2176 1469
rect 2182 1463 2186 1469
rect 2206 1463 2210 1469
rect 2214 1463 2218 1469
rect 2253 1463 2257 1469
rect 2262 1463 2266 1469
rect 2272 1463 2276 1469
rect 2296 1463 2300 1469
rect 2304 1463 2308 1469
rect 2348 1463 2352 1469
rect 2357 1463 2361 1469
rect 2367 1463 2371 1469
rect 2391 1463 2395 1469
rect 2399 1463 2403 1469
rect 3481 1469 3485 1475
rect 3490 1469 3494 1475
rect 3500 1469 3504 1475
rect 3510 1469 3514 1475
rect 3520 1469 3524 1475
rect 3542 1469 3546 1475
rect 3550 1469 3554 1475
rect 3024 1455 3028 1461
rect 3033 1455 3037 1461
rect 3043 1455 3047 1461
rect 3067 1455 3071 1461
rect 3075 1455 3079 1461
rect 3226 1460 3230 1466
rect 3235 1460 3239 1466
rect 3245 1460 3249 1466
rect 3255 1460 3259 1466
rect 3279 1460 3283 1466
rect 3287 1460 3291 1466
rect 4003 1408 4007 1414
rect 4041 1408 4045 1414
rect 4051 1408 4055 1414
rect 4059 1408 4063 1414
rect 1012 1389 1016 1395
rect 1021 1389 1025 1395
rect 1031 1389 1035 1395
rect 1055 1389 1059 1395
rect 1063 1389 1067 1395
rect 3084 1294 3088 1298
rect 3092 1294 3096 1298
rect 3140 1294 3144 1298
rect 3148 1294 3152 1298
rect 3337 1294 3341 1298
rect 3345 1294 3349 1298
rect 3600 1294 3604 1298
rect 3608 1294 3612 1298
rect 1766 1146 1770 1152
rect 1775 1146 1779 1152
rect 1785 1146 1789 1152
rect 1809 1146 1813 1152
rect 1817 1146 1821 1152
rect 1852 1146 1856 1152
rect 1861 1146 1865 1152
rect 1871 1146 1875 1152
rect 1895 1146 1899 1152
rect 1903 1146 1907 1152
rect 1942 1146 1946 1152
rect 1951 1146 1955 1152
rect 1961 1146 1965 1152
rect 1985 1146 1989 1152
rect 1993 1146 1997 1152
rect 2037 1146 2041 1152
rect 2046 1146 2050 1152
rect 2056 1146 2060 1152
rect 2080 1146 2084 1152
rect 2088 1146 2092 1152
rect 2121 1146 2125 1152
rect 2130 1146 2134 1152
rect 2140 1146 2144 1152
rect 2164 1146 2168 1152
rect 2172 1146 2176 1152
rect 2207 1146 2211 1152
rect 2216 1146 2220 1152
rect 2226 1146 2230 1152
rect 2250 1146 2254 1152
rect 2258 1146 2262 1152
rect 2297 1146 2301 1152
rect 2306 1146 2310 1152
rect 2316 1146 2320 1152
rect 2340 1146 2344 1152
rect 2348 1146 2352 1152
rect 2392 1146 2396 1152
rect 2401 1146 2405 1152
rect 2411 1146 2415 1152
rect 2435 1146 2439 1152
rect 2443 1146 2447 1152
rect 1828 1045 1832 1051
rect 1837 1045 1841 1051
rect 1847 1045 1851 1051
rect 1871 1045 1875 1051
rect 1879 1045 1883 1051
rect 1914 1045 1918 1051
rect 1923 1045 1927 1051
rect 1933 1045 1937 1051
rect 1957 1045 1961 1051
rect 1965 1045 1969 1051
rect 2004 1045 2008 1051
rect 2013 1045 2017 1051
rect 2023 1045 2027 1051
rect 2047 1045 2051 1051
rect 2055 1045 2059 1051
rect 2099 1045 2103 1051
rect 2108 1045 2112 1051
rect 2118 1045 2122 1051
rect 2142 1045 2146 1051
rect 2150 1045 2154 1051
<< polysilicon >>
rect 2015 3429 2101 3431
rect 2015 3421 2017 3429
rect 2031 3421 2033 3424
rect 2041 3421 2043 3424
rect 2051 3421 2053 3429
rect 2061 3421 2063 3424
rect 2081 3421 2083 3424
rect 1778 3419 1864 3421
rect 1616 3410 1702 3412
rect 1778 3411 1780 3419
rect 1794 3411 1796 3414
rect 1804 3411 1806 3414
rect 1814 3411 1816 3419
rect 1824 3411 1826 3414
rect 1844 3411 1846 3414
rect 1616 3402 1618 3410
rect 1632 3402 1634 3405
rect 1642 3402 1644 3405
rect 1652 3402 1654 3410
rect 1662 3402 1664 3405
rect 1682 3402 1684 3405
rect 1616 3354 1618 3396
rect 1632 3354 1634 3396
rect 1642 3375 1644 3396
rect 1652 3393 1654 3396
rect 1642 3373 1654 3375
rect 1642 3354 1644 3357
rect 1652 3354 1654 3373
rect 1662 3354 1664 3396
rect 1682 3373 1684 3396
rect 1700 3368 1702 3410
rect 1673 3366 1702 3368
rect 1616 3347 1618 3350
rect 1632 3339 1634 3350
rect 1642 3344 1644 3350
rect 1652 3347 1654 3350
rect 1662 3347 1664 3350
rect 1673 3344 1675 3366
rect 1778 3363 1780 3405
rect 1794 3363 1796 3405
rect 1804 3384 1806 3405
rect 1814 3402 1816 3405
rect 1804 3382 1816 3384
rect 1804 3363 1806 3366
rect 1814 3363 1816 3382
rect 1824 3363 1826 3405
rect 1844 3382 1846 3405
rect 1862 3377 1864 3419
rect 1835 3375 1864 3377
rect 1682 3354 1684 3362
rect 1778 3356 1780 3359
rect 1642 3342 1675 3344
rect 1682 3339 1684 3350
rect 1794 3348 1796 3359
rect 1804 3353 1806 3359
rect 1814 3356 1816 3359
rect 1824 3356 1826 3359
rect 1835 3353 1837 3375
rect 2015 3373 2017 3415
rect 2031 3373 2033 3415
rect 2041 3394 2043 3415
rect 2051 3412 2053 3415
rect 2041 3392 2053 3394
rect 2041 3373 2043 3376
rect 2051 3373 2053 3392
rect 2061 3373 2063 3415
rect 2081 3392 2083 3415
rect 2099 3387 2101 3429
rect 2072 3385 2101 3387
rect 1844 3363 1846 3371
rect 2015 3366 2017 3369
rect 1804 3351 1837 3353
rect 1844 3348 1846 3359
rect 2031 3358 2033 3369
rect 2041 3363 2043 3369
rect 2051 3366 2053 3369
rect 2061 3366 2063 3369
rect 2072 3363 2074 3385
rect 2081 3373 2083 3381
rect 2041 3361 2074 3363
rect 2081 3358 2083 3369
rect 2031 3356 2083 3358
rect 1794 3346 1846 3348
rect 1632 3337 1684 3339
rect 1904 3295 1906 3304
rect 1914 3295 1916 3304
rect 1947 3295 1949 3304
rect 2032 3296 2034 3305
rect 2042 3296 2044 3305
rect 2075 3296 2077 3305
rect 1904 3263 1906 3289
rect 1914 3263 1916 3289
rect 1947 3263 1949 3289
rect 2032 3264 2034 3290
rect 2042 3264 2044 3290
rect 2075 3264 2077 3290
rect 1904 3256 1906 3259
rect 1914 3256 1916 3259
rect 1947 3256 1949 3259
rect 2032 3257 2034 3260
rect 2042 3257 2044 3260
rect 2075 3257 2077 3260
rect 2073 3224 2075 3227
rect 2083 3224 2085 3227
rect 2101 3224 2103 3227
rect 2073 3186 2075 3218
rect 2083 3186 2085 3218
rect 2101 3186 2103 3218
rect 2073 3179 2075 3182
rect 2083 3179 2085 3182
rect 2101 3179 2103 3182
rect 2024 3097 2110 3099
rect 2024 3089 2026 3097
rect 2040 3089 2042 3092
rect 2050 3089 2052 3092
rect 2060 3089 2062 3097
rect 2070 3089 2072 3092
rect 2090 3089 2092 3092
rect 1787 3087 1873 3089
rect 1625 3078 1711 3080
rect 1787 3079 1789 3087
rect 1803 3079 1805 3082
rect 1813 3079 1815 3082
rect 1823 3079 1825 3087
rect 1833 3079 1835 3082
rect 1853 3079 1855 3082
rect 1625 3070 1627 3078
rect 1641 3070 1643 3073
rect 1651 3070 1653 3073
rect 1661 3070 1663 3078
rect 1671 3070 1673 3073
rect 1691 3070 1693 3073
rect 1625 3022 1627 3064
rect 1641 3022 1643 3064
rect 1651 3043 1653 3064
rect 1661 3061 1663 3064
rect 1651 3041 1663 3043
rect 1651 3022 1653 3025
rect 1661 3022 1663 3041
rect 1671 3022 1673 3064
rect 1691 3041 1693 3064
rect 1709 3036 1711 3078
rect 1682 3034 1711 3036
rect 1625 3015 1627 3018
rect 1641 3007 1643 3018
rect 1651 3012 1653 3018
rect 1661 3015 1663 3018
rect 1671 3015 1673 3018
rect 1682 3012 1684 3034
rect 1787 3031 1789 3073
rect 1803 3031 1805 3073
rect 1813 3052 1815 3073
rect 1823 3070 1825 3073
rect 1813 3050 1825 3052
rect 1813 3031 1815 3034
rect 1823 3031 1825 3050
rect 1833 3031 1835 3073
rect 1853 3050 1855 3073
rect 1871 3045 1873 3087
rect 1844 3043 1873 3045
rect 1691 3022 1693 3030
rect 1787 3024 1789 3027
rect 1651 3010 1684 3012
rect 1691 3007 1693 3018
rect 1803 3016 1805 3027
rect 1813 3021 1815 3027
rect 1823 3024 1825 3027
rect 1833 3024 1835 3027
rect 1844 3021 1846 3043
rect 2024 3041 2026 3083
rect 2040 3041 2042 3083
rect 2050 3062 2052 3083
rect 2060 3080 2062 3083
rect 2050 3060 2062 3062
rect 2050 3041 2052 3044
rect 2060 3041 2062 3060
rect 2070 3041 2072 3083
rect 2090 3060 2092 3083
rect 2108 3055 2110 3097
rect 2081 3053 2110 3055
rect 1853 3031 1855 3039
rect 2024 3034 2026 3037
rect 1813 3019 1846 3021
rect 1853 3016 1855 3027
rect 2040 3026 2042 3037
rect 2050 3031 2052 3037
rect 2060 3034 2062 3037
rect 2070 3034 2072 3037
rect 2081 3031 2083 3053
rect 2090 3041 2092 3049
rect 2050 3029 2083 3031
rect 2090 3026 2092 3037
rect 2040 3024 2092 3026
rect 1803 3014 1855 3016
rect 1641 3005 1693 3007
rect 1913 2963 1915 2972
rect 1923 2963 1925 2972
rect 1956 2963 1958 2972
rect 2041 2964 2043 2973
rect 2051 2964 2053 2973
rect 2084 2964 2086 2973
rect 1913 2931 1915 2957
rect 1923 2931 1925 2957
rect 1956 2931 1958 2957
rect 2041 2932 2043 2958
rect 2051 2932 2053 2958
rect 2084 2932 2086 2958
rect 1913 2924 1915 2927
rect 1923 2924 1925 2927
rect 1956 2924 1958 2927
rect 2041 2925 2043 2928
rect 2051 2925 2053 2928
rect 2084 2925 2086 2928
rect 2082 2892 2084 2895
rect 2092 2892 2094 2895
rect 2110 2892 2112 2895
rect 2082 2854 2084 2886
rect 2092 2854 2094 2886
rect 2110 2854 2112 2886
rect 2082 2847 2084 2850
rect 2092 2847 2094 2850
rect 2110 2847 2112 2850
rect 2045 2731 2131 2733
rect 2045 2723 2047 2731
rect 2061 2723 2063 2726
rect 2071 2723 2073 2726
rect 2081 2723 2083 2731
rect 2091 2723 2093 2726
rect 2111 2723 2113 2726
rect 1808 2721 1894 2723
rect 1646 2712 1732 2714
rect 1808 2713 1810 2721
rect 1824 2713 1826 2716
rect 1834 2713 1836 2716
rect 1844 2713 1846 2721
rect 1854 2713 1856 2716
rect 1874 2713 1876 2716
rect 1646 2704 1648 2712
rect 1662 2704 1664 2707
rect 1672 2704 1674 2707
rect 1682 2704 1684 2712
rect 1692 2704 1694 2707
rect 1712 2704 1714 2707
rect 1646 2656 1648 2698
rect 1662 2656 1664 2698
rect 1672 2677 1674 2698
rect 1682 2695 1684 2698
rect 1672 2675 1684 2677
rect 1672 2656 1674 2659
rect 1682 2656 1684 2675
rect 1692 2656 1694 2698
rect 1712 2675 1714 2698
rect 1730 2670 1732 2712
rect 1703 2668 1732 2670
rect 1646 2649 1648 2652
rect 1662 2641 1664 2652
rect 1672 2646 1674 2652
rect 1682 2649 1684 2652
rect 1692 2649 1694 2652
rect 1703 2646 1705 2668
rect 1808 2665 1810 2707
rect 1824 2665 1826 2707
rect 1834 2686 1836 2707
rect 1844 2704 1846 2707
rect 1834 2684 1846 2686
rect 1834 2665 1836 2668
rect 1844 2665 1846 2684
rect 1854 2665 1856 2707
rect 1874 2684 1876 2707
rect 1892 2679 1894 2721
rect 1865 2677 1894 2679
rect 1712 2656 1714 2664
rect 1808 2658 1810 2661
rect 1672 2644 1705 2646
rect 1712 2641 1714 2652
rect 1824 2650 1826 2661
rect 1834 2655 1836 2661
rect 1844 2658 1846 2661
rect 1854 2658 1856 2661
rect 1865 2655 1867 2677
rect 2045 2675 2047 2717
rect 2061 2675 2063 2717
rect 2071 2696 2073 2717
rect 2081 2714 2083 2717
rect 2071 2694 2083 2696
rect 2071 2675 2073 2678
rect 2081 2675 2083 2694
rect 2091 2675 2093 2717
rect 2111 2694 2113 2717
rect 2129 2689 2131 2731
rect 2102 2687 2131 2689
rect 1874 2665 1876 2673
rect 2045 2668 2047 2671
rect 1834 2653 1867 2655
rect 1874 2650 1876 2661
rect 2061 2660 2063 2671
rect 2071 2665 2073 2671
rect 2081 2668 2083 2671
rect 2091 2668 2093 2671
rect 2102 2665 2104 2687
rect 2111 2675 2113 2683
rect 2071 2663 2104 2665
rect 2111 2660 2113 2671
rect 2061 2658 2113 2660
rect 1824 2648 1876 2650
rect 1662 2639 1714 2641
rect 1934 2597 1936 2606
rect 1944 2597 1946 2606
rect 1977 2597 1979 2606
rect 2062 2598 2064 2607
rect 2072 2598 2074 2607
rect 2105 2598 2107 2607
rect 1934 2565 1936 2591
rect 1944 2565 1946 2591
rect 1977 2565 1979 2591
rect 2062 2566 2064 2592
rect 2072 2566 2074 2592
rect 2105 2566 2107 2592
rect 1934 2558 1936 2561
rect 1944 2558 1946 2561
rect 1977 2558 1979 2561
rect 2062 2559 2064 2562
rect 2072 2559 2074 2562
rect 2105 2559 2107 2562
rect 2103 2526 2105 2529
rect 2113 2526 2115 2529
rect 2131 2526 2133 2529
rect 2103 2488 2105 2520
rect 2113 2488 2115 2520
rect 2131 2488 2133 2520
rect 2103 2481 2105 2484
rect 2113 2481 2115 2484
rect 2131 2481 2133 2484
rect 2073 2357 2159 2359
rect 2073 2349 2075 2357
rect 2089 2349 2091 2352
rect 2099 2349 2101 2352
rect 2109 2349 2111 2357
rect 2119 2349 2121 2352
rect 2139 2349 2141 2352
rect 1836 2347 1922 2349
rect 1674 2338 1760 2340
rect 1836 2339 1838 2347
rect 1852 2339 1854 2342
rect 1862 2339 1864 2342
rect 1872 2339 1874 2347
rect 1882 2339 1884 2342
rect 1902 2339 1904 2342
rect 1674 2330 1676 2338
rect 1690 2330 1692 2333
rect 1700 2330 1702 2333
rect 1710 2330 1712 2338
rect 1720 2330 1722 2333
rect 1740 2330 1742 2333
rect 1674 2282 1676 2324
rect 1690 2282 1692 2324
rect 1700 2303 1702 2324
rect 1710 2321 1712 2324
rect 1700 2301 1712 2303
rect 1700 2282 1702 2285
rect 1710 2282 1712 2301
rect 1720 2282 1722 2324
rect 1740 2301 1742 2324
rect 1758 2296 1760 2338
rect 1731 2294 1760 2296
rect 1674 2275 1676 2278
rect 1690 2267 1692 2278
rect 1700 2272 1702 2278
rect 1710 2275 1712 2278
rect 1720 2275 1722 2278
rect 1731 2272 1733 2294
rect 1836 2291 1838 2333
rect 1852 2291 1854 2333
rect 1862 2312 1864 2333
rect 1872 2330 1874 2333
rect 1862 2310 1874 2312
rect 1862 2291 1864 2294
rect 1872 2291 1874 2310
rect 1882 2291 1884 2333
rect 1902 2310 1904 2333
rect 1920 2305 1922 2347
rect 1893 2303 1922 2305
rect 1740 2282 1742 2290
rect 1836 2284 1838 2287
rect 1700 2270 1733 2272
rect 1740 2267 1742 2278
rect 1852 2276 1854 2287
rect 1862 2281 1864 2287
rect 1872 2284 1874 2287
rect 1882 2284 1884 2287
rect 1893 2281 1895 2303
rect 2073 2301 2075 2343
rect 2089 2301 2091 2343
rect 2099 2322 2101 2343
rect 2109 2340 2111 2343
rect 2099 2320 2111 2322
rect 2099 2301 2101 2304
rect 2109 2301 2111 2320
rect 2119 2301 2121 2343
rect 2139 2320 2141 2343
rect 2157 2315 2159 2357
rect 2130 2313 2159 2315
rect 1902 2291 1904 2299
rect 2073 2294 2075 2297
rect 1862 2279 1895 2281
rect 1902 2276 1904 2287
rect 2089 2286 2091 2297
rect 2099 2291 2101 2297
rect 2109 2294 2111 2297
rect 2119 2294 2121 2297
rect 2130 2291 2132 2313
rect 2139 2301 2141 2309
rect 2099 2289 2132 2291
rect 2139 2286 2141 2297
rect 2089 2284 2141 2286
rect 1852 2274 1904 2276
rect 1690 2265 1742 2267
rect 1962 2223 1964 2232
rect 1972 2223 1974 2232
rect 2005 2223 2007 2232
rect 2090 2224 2092 2233
rect 2100 2224 2102 2233
rect 2133 2224 2135 2233
rect 1962 2191 1964 2217
rect 1972 2191 1974 2217
rect 2005 2191 2007 2217
rect 2090 2192 2092 2218
rect 2100 2192 2102 2218
rect 2133 2192 2135 2218
rect 1962 2184 1964 2187
rect 1972 2184 1974 2187
rect 2005 2184 2007 2187
rect 2090 2185 2092 2188
rect 2100 2185 2102 2188
rect 2133 2185 2135 2188
rect 2131 2152 2133 2155
rect 2141 2152 2143 2155
rect 2159 2152 2161 2155
rect 2131 2114 2133 2146
rect 2141 2114 2143 2146
rect 2159 2114 2161 2146
rect 2131 2107 2133 2110
rect 2141 2107 2143 2110
rect 2159 2107 2161 2110
rect 3959 1787 3961 1796
rect 3969 1787 3971 1796
rect 3979 1787 3981 1796
rect 3989 1787 3991 1796
rect 4020 1787 4022 1796
rect 3959 1744 3961 1781
rect 3969 1744 3971 1781
rect 3979 1744 3981 1781
rect 3989 1744 3991 1781
rect 4020 1744 4022 1781
rect 3959 1737 3961 1740
rect 3969 1737 3971 1740
rect 3979 1737 3981 1740
rect 3989 1737 3991 1740
rect 4020 1737 4022 1740
rect 1053 1727 1055 1730
rect 1109 1727 1111 1730
rect 1053 1714 1055 1723
rect 1049 1712 1055 1714
rect 1053 1707 1055 1712
rect 1109 1714 1111 1723
rect 1105 1712 1111 1714
rect 1749 1713 1751 1722
rect 1759 1713 1761 1722
rect 1792 1713 1794 1722
rect 1835 1713 1837 1722
rect 1845 1713 1847 1722
rect 1878 1713 1880 1722
rect 1925 1713 1927 1722
rect 1935 1713 1937 1722
rect 1968 1713 1970 1722
rect 2020 1713 2022 1722
rect 2030 1713 2032 1722
rect 2063 1713 2065 1722
rect 2104 1713 2106 1722
rect 2114 1713 2116 1722
rect 2147 1713 2149 1722
rect 2190 1713 2192 1722
rect 2200 1713 2202 1722
rect 2233 1713 2235 1722
rect 2280 1713 2282 1722
rect 2290 1713 2292 1722
rect 2323 1713 2325 1722
rect 2375 1713 2377 1722
rect 2385 1713 2387 1722
rect 2418 1713 2420 1722
rect 1109 1707 1111 1712
rect 1053 1700 1055 1703
rect 1109 1700 1111 1703
rect 1749 1681 1751 1707
rect 1759 1681 1761 1707
rect 1792 1681 1794 1707
rect 1835 1681 1837 1707
rect 1845 1681 1847 1707
rect 1878 1681 1880 1707
rect 1925 1681 1927 1707
rect 1935 1681 1937 1707
rect 1968 1681 1970 1707
rect 2020 1681 2022 1707
rect 2030 1681 2032 1707
rect 2063 1681 2065 1707
rect 2104 1681 2106 1707
rect 2114 1681 2116 1707
rect 2147 1681 2149 1707
rect 2190 1681 2192 1707
rect 2200 1681 2202 1707
rect 2233 1681 2235 1707
rect 2280 1681 2282 1707
rect 2290 1681 2292 1707
rect 2323 1681 2325 1707
rect 2375 1681 2377 1707
rect 2385 1681 2387 1707
rect 2418 1681 2420 1707
rect 1749 1674 1751 1677
rect 1759 1674 1761 1677
rect 1792 1674 1794 1677
rect 1835 1674 1837 1677
rect 1845 1674 1847 1677
rect 1878 1674 1880 1677
rect 1925 1674 1927 1677
rect 1935 1674 1937 1677
rect 1968 1674 1970 1677
rect 2020 1674 2022 1677
rect 2030 1674 2032 1677
rect 2063 1674 2065 1677
rect 2104 1674 2106 1677
rect 2114 1674 2116 1677
rect 2147 1674 2149 1677
rect 2190 1674 2192 1677
rect 2200 1674 2202 1677
rect 2233 1674 2235 1677
rect 2280 1674 2282 1677
rect 2290 1674 2292 1677
rect 2323 1674 2325 1677
rect 2375 1674 2377 1677
rect 2385 1674 2387 1677
rect 2418 1674 2420 1677
rect 2964 1669 3050 1671
rect 2964 1661 2966 1669
rect 2980 1661 2982 1664
rect 2990 1661 2992 1664
rect 3000 1661 3002 1669
rect 3010 1661 3012 1664
rect 3030 1661 3032 1664
rect 1016 1652 1018 1661
rect 1026 1652 1028 1661
rect 1059 1652 1061 1661
rect 1016 1620 1018 1646
rect 1026 1620 1028 1646
rect 1059 1620 1061 1646
rect 1016 1613 1018 1616
rect 1026 1613 1028 1616
rect 1059 1613 1061 1616
rect 2964 1613 2966 1655
rect 2980 1613 2982 1655
rect 2990 1634 2992 1655
rect 3000 1652 3002 1655
rect 2990 1632 3002 1634
rect 2990 1613 2992 1616
rect 3000 1613 3002 1632
rect 3010 1613 3012 1655
rect 3030 1632 3032 1655
rect 3048 1627 3050 1669
rect 3213 1669 3299 1671
rect 3213 1661 3215 1669
rect 3229 1661 3231 1664
rect 3239 1661 3241 1664
rect 3249 1661 3251 1669
rect 3259 1661 3261 1664
rect 3279 1661 3281 1664
rect 3104 1656 3106 1659
rect 3104 1643 3106 1652
rect 3100 1641 3106 1643
rect 3104 1636 3106 1641
rect 3104 1629 3106 1632
rect 3021 1625 3050 1627
rect 2964 1606 2966 1609
rect 2980 1598 2982 1609
rect 2990 1603 2992 1609
rect 3000 1606 3002 1609
rect 3010 1606 3012 1609
rect 3021 1603 3023 1625
rect 3030 1613 3032 1621
rect 3213 1613 3215 1655
rect 3229 1613 3231 1655
rect 3239 1634 3241 1655
rect 3249 1652 3251 1655
rect 3239 1632 3251 1634
rect 3239 1613 3241 1616
rect 3249 1613 3251 1632
rect 3259 1613 3261 1655
rect 3279 1632 3281 1655
rect 3297 1627 3299 1669
rect 3470 1669 3556 1671
rect 3470 1661 3472 1669
rect 3486 1661 3488 1664
rect 3496 1661 3498 1664
rect 3506 1661 3508 1669
rect 3516 1661 3518 1664
rect 3536 1661 3538 1664
rect 3353 1656 3355 1659
rect 3353 1643 3355 1652
rect 3349 1641 3355 1643
rect 3353 1636 3355 1641
rect 3353 1629 3355 1632
rect 3270 1625 3299 1627
rect 2990 1601 3023 1603
rect 3030 1598 3032 1609
rect 3213 1606 3215 1609
rect 2980 1596 3032 1598
rect 3229 1598 3231 1609
rect 3239 1603 3241 1609
rect 3249 1606 3251 1609
rect 3259 1606 3261 1609
rect 3270 1603 3272 1625
rect 3279 1613 3281 1621
rect 3470 1613 3472 1655
rect 3486 1613 3488 1655
rect 3496 1634 3498 1655
rect 3506 1652 3508 1655
rect 3496 1632 3508 1634
rect 3496 1613 3498 1616
rect 3506 1613 3508 1632
rect 3516 1613 3518 1655
rect 3536 1632 3538 1655
rect 3554 1627 3556 1669
rect 3692 1669 3778 1671
rect 3692 1661 3694 1669
rect 3708 1661 3710 1664
rect 3718 1661 3720 1664
rect 3728 1661 3730 1669
rect 3738 1661 3740 1664
rect 3758 1661 3760 1664
rect 3610 1656 3612 1659
rect 3610 1643 3612 1652
rect 3606 1641 3612 1643
rect 3610 1636 3612 1641
rect 3610 1629 3612 1632
rect 3527 1625 3556 1627
rect 3239 1601 3272 1603
rect 3279 1598 3281 1609
rect 3470 1606 3472 1609
rect 3229 1596 3281 1598
rect 3486 1598 3488 1609
rect 3496 1603 3498 1609
rect 3506 1606 3508 1609
rect 3516 1606 3518 1609
rect 3527 1603 3529 1625
rect 3536 1613 3538 1621
rect 3692 1613 3694 1655
rect 3708 1613 3710 1655
rect 3718 1634 3720 1655
rect 3728 1652 3730 1655
rect 3718 1632 3730 1634
rect 3718 1613 3720 1616
rect 3728 1613 3730 1632
rect 3738 1613 3740 1655
rect 3758 1632 3760 1655
rect 3776 1627 3778 1669
rect 3832 1656 3834 1659
rect 3832 1643 3834 1652
rect 3828 1641 3834 1643
rect 3832 1636 3834 1641
rect 4258 1632 4260 1635
rect 4268 1632 4270 1635
rect 3832 1629 3834 1632
rect 3749 1625 3778 1627
rect 3496 1601 3529 1603
rect 3536 1598 3538 1609
rect 3692 1606 3694 1609
rect 3486 1596 3538 1598
rect 3708 1598 3710 1609
rect 3718 1603 3720 1609
rect 3728 1606 3730 1609
rect 3738 1606 3740 1609
rect 3749 1603 3751 1625
rect 3758 1613 3760 1621
rect 3718 1601 3751 1603
rect 3758 1598 3760 1609
rect 3708 1596 3760 1598
rect 4258 1594 4260 1626
rect 4268 1594 4270 1626
rect 4258 1587 4260 1590
rect 4268 1587 4270 1590
rect 1322 1581 1324 1584
rect 1332 1581 1334 1584
rect 1350 1581 1352 1584
rect 1017 1567 1019 1576
rect 1027 1567 1029 1576
rect 1060 1567 1062 1576
rect 1017 1535 1019 1561
rect 1027 1535 1029 1561
rect 1060 1535 1062 1561
rect 1322 1543 1324 1575
rect 1332 1543 1334 1575
rect 1350 1543 1352 1575
rect 1322 1536 1324 1539
rect 1332 1536 1334 1539
rect 1350 1536 1352 1539
rect 1017 1528 1019 1531
rect 1027 1528 1029 1531
rect 1060 1528 1062 1531
rect 1017 1478 1019 1487
rect 1027 1478 1029 1487
rect 1060 1478 1062 1487
rect 3747 1485 3749 1494
rect 3757 1485 3759 1494
rect 3767 1485 3769 1494
rect 3777 1485 3779 1494
rect 3787 1485 3789 1494
rect 3820 1485 3822 1494
rect 1017 1446 1019 1472
rect 1027 1446 1029 1472
rect 1060 1446 1062 1472
rect 1727 1469 1729 1478
rect 1737 1469 1739 1478
rect 1770 1469 1772 1478
rect 1813 1469 1815 1478
rect 1823 1469 1825 1478
rect 1856 1469 1858 1478
rect 1903 1469 1905 1478
rect 1913 1469 1915 1478
rect 1946 1469 1948 1478
rect 1998 1469 2000 1478
rect 2008 1469 2010 1478
rect 2041 1469 2043 1478
rect 2082 1469 2084 1478
rect 2092 1469 2094 1478
rect 2125 1469 2127 1478
rect 2168 1469 2170 1478
rect 2178 1469 2180 1478
rect 2211 1469 2213 1478
rect 2258 1469 2260 1478
rect 2268 1469 2270 1478
rect 2301 1469 2303 1478
rect 2353 1469 2355 1478
rect 2363 1469 2365 1478
rect 2396 1469 2398 1478
rect 3486 1475 3488 1484
rect 3496 1475 3498 1484
rect 3506 1475 3508 1484
rect 3516 1475 3518 1484
rect 3547 1475 3549 1484
rect 1017 1439 1019 1442
rect 1027 1439 1029 1442
rect 1060 1439 1062 1442
rect 1727 1437 1729 1463
rect 1737 1437 1739 1463
rect 1770 1437 1772 1463
rect 1813 1437 1815 1463
rect 1823 1437 1825 1463
rect 1856 1437 1858 1463
rect 1903 1437 1905 1463
rect 1913 1437 1915 1463
rect 1946 1437 1948 1463
rect 1998 1437 2000 1463
rect 2008 1437 2010 1463
rect 2041 1437 2043 1463
rect 2082 1437 2084 1463
rect 2092 1437 2094 1463
rect 2125 1437 2127 1463
rect 2168 1437 2170 1463
rect 2178 1437 2180 1463
rect 2211 1437 2213 1463
rect 2258 1437 2260 1463
rect 2268 1437 2270 1463
rect 2301 1437 2303 1463
rect 2353 1437 2355 1463
rect 2363 1437 2365 1463
rect 2396 1437 2398 1463
rect 3029 1461 3031 1470
rect 3039 1461 3041 1470
rect 3072 1461 3074 1470
rect 3231 1466 3233 1475
rect 3241 1466 3243 1475
rect 3251 1466 3253 1475
rect 3284 1466 3286 1475
rect 1727 1430 1729 1433
rect 1737 1430 1739 1433
rect 1770 1430 1772 1433
rect 1813 1430 1815 1433
rect 1823 1430 1825 1433
rect 1856 1430 1858 1433
rect 1903 1430 1905 1433
rect 1913 1430 1915 1433
rect 1946 1430 1948 1433
rect 1998 1430 2000 1433
rect 2008 1430 2010 1433
rect 2041 1430 2043 1433
rect 2082 1430 2084 1433
rect 2092 1430 2094 1433
rect 2125 1430 2127 1433
rect 2168 1430 2170 1433
rect 2178 1430 2180 1433
rect 2211 1430 2213 1433
rect 2258 1430 2260 1433
rect 2268 1430 2270 1433
rect 2301 1430 2303 1433
rect 2353 1430 2355 1433
rect 2363 1430 2365 1433
rect 2396 1430 2398 1433
rect 3029 1429 3031 1455
rect 3039 1429 3041 1455
rect 3072 1429 3074 1455
rect 3231 1431 3233 1460
rect 3241 1431 3243 1460
rect 3251 1431 3253 1460
rect 3284 1431 3286 1460
rect 3486 1432 3488 1469
rect 3496 1432 3498 1469
rect 3506 1432 3508 1469
rect 3516 1432 3518 1469
rect 3547 1432 3549 1469
rect 3747 1435 3749 1479
rect 3757 1435 3759 1479
rect 3767 1435 3769 1479
rect 3777 1435 3779 1479
rect 3787 1435 3789 1479
rect 3820 1435 3822 1479
rect 3747 1428 3749 1431
rect 3757 1428 3759 1431
rect 3767 1428 3769 1431
rect 3777 1428 3779 1431
rect 3787 1428 3789 1431
rect 3820 1428 3822 1431
rect 3029 1422 3031 1425
rect 3039 1422 3041 1425
rect 3072 1422 3074 1425
rect 3231 1424 3233 1427
rect 3241 1424 3243 1427
rect 3251 1424 3253 1427
rect 3284 1424 3286 1427
rect 3486 1425 3488 1428
rect 3496 1425 3498 1428
rect 3506 1425 3508 1428
rect 3516 1425 3518 1428
rect 3547 1425 3549 1428
rect 4008 1414 4010 1417
rect 4018 1414 4020 1417
rect 4027 1414 4029 1417
rect 4037 1414 4039 1417
rect 4056 1414 4058 1417
rect 1017 1395 1019 1404
rect 1027 1395 1029 1404
rect 1060 1395 1062 1404
rect 1017 1363 1019 1389
rect 1027 1363 1029 1389
rect 1060 1363 1062 1389
rect 4008 1362 4010 1408
rect 4018 1362 4020 1408
rect 4027 1385 4029 1408
rect 4028 1381 4029 1385
rect 4027 1362 4029 1381
rect 4037 1362 4039 1408
rect 4056 1362 4058 1408
rect 1017 1356 1019 1359
rect 1027 1356 1029 1359
rect 1060 1356 1062 1359
rect 4008 1355 4010 1358
rect 4018 1355 4020 1358
rect 4027 1355 4029 1358
rect 4037 1355 4039 1358
rect 4056 1355 4058 1358
rect 3089 1298 3091 1301
rect 3145 1298 3147 1301
rect 3342 1298 3344 1301
rect 3605 1298 3607 1301
rect 3089 1285 3091 1294
rect 3085 1283 3091 1285
rect 3089 1278 3091 1283
rect 3145 1285 3147 1294
rect 3141 1283 3147 1285
rect 3145 1278 3147 1283
rect 3342 1285 3344 1294
rect 3338 1283 3344 1285
rect 3342 1278 3344 1283
rect 3605 1285 3607 1294
rect 3601 1283 3607 1285
rect 3605 1278 3607 1283
rect 3089 1271 3091 1274
rect 3145 1271 3147 1274
rect 3342 1271 3344 1274
rect 3605 1271 3607 1274
rect 1771 1152 1773 1161
rect 1781 1152 1783 1161
rect 1814 1152 1816 1161
rect 1857 1152 1859 1161
rect 1867 1152 1869 1161
rect 1900 1152 1902 1161
rect 1947 1152 1949 1161
rect 1957 1152 1959 1161
rect 1990 1152 1992 1161
rect 2042 1152 2044 1161
rect 2052 1152 2054 1161
rect 2085 1152 2087 1161
rect 2126 1152 2128 1161
rect 2136 1152 2138 1161
rect 2169 1152 2171 1161
rect 2212 1152 2214 1161
rect 2222 1152 2224 1161
rect 2255 1152 2257 1161
rect 2302 1152 2304 1161
rect 2312 1152 2314 1161
rect 2345 1152 2347 1161
rect 2397 1152 2399 1161
rect 2407 1152 2409 1161
rect 2440 1152 2442 1161
rect 1771 1120 1773 1146
rect 1781 1120 1783 1146
rect 1814 1120 1816 1146
rect 1857 1120 1859 1146
rect 1867 1120 1869 1146
rect 1900 1120 1902 1146
rect 1947 1120 1949 1146
rect 1957 1120 1959 1146
rect 1990 1120 1992 1146
rect 2042 1120 2044 1146
rect 2052 1120 2054 1146
rect 2085 1120 2087 1146
rect 2126 1120 2128 1146
rect 2136 1120 2138 1146
rect 2169 1120 2171 1146
rect 2212 1120 2214 1146
rect 2222 1120 2224 1146
rect 2255 1120 2257 1146
rect 2302 1120 2304 1146
rect 2312 1120 2314 1146
rect 2345 1120 2347 1146
rect 2397 1120 2399 1146
rect 2407 1120 2409 1146
rect 2440 1120 2442 1146
rect 1771 1113 1773 1116
rect 1781 1113 1783 1116
rect 1814 1113 1816 1116
rect 1857 1113 1859 1116
rect 1867 1113 1869 1116
rect 1900 1113 1902 1116
rect 1947 1113 1949 1116
rect 1957 1113 1959 1116
rect 1990 1113 1992 1116
rect 2042 1113 2044 1116
rect 2052 1113 2054 1116
rect 2085 1113 2087 1116
rect 2126 1113 2128 1116
rect 2136 1113 2138 1116
rect 2169 1113 2171 1116
rect 2212 1113 2214 1116
rect 2222 1113 2224 1116
rect 2255 1113 2257 1116
rect 2302 1113 2304 1116
rect 2312 1113 2314 1116
rect 2345 1113 2347 1116
rect 2397 1113 2399 1116
rect 2407 1113 2409 1116
rect 2440 1113 2442 1116
rect 1833 1051 1835 1060
rect 1843 1051 1845 1060
rect 1876 1051 1878 1060
rect 1919 1051 1921 1060
rect 1929 1051 1931 1060
rect 1962 1051 1964 1060
rect 2009 1051 2011 1060
rect 2019 1051 2021 1060
rect 2052 1051 2054 1060
rect 2104 1051 2106 1060
rect 2114 1051 2116 1060
rect 2147 1051 2149 1060
rect 1833 1019 1835 1045
rect 1843 1019 1845 1045
rect 1876 1019 1878 1045
rect 1919 1019 1921 1045
rect 1929 1019 1931 1045
rect 1962 1019 1964 1045
rect 2009 1019 2011 1045
rect 2019 1019 2021 1045
rect 2052 1019 2054 1045
rect 2104 1019 2106 1045
rect 2114 1019 2116 1045
rect 2147 1019 2149 1045
rect 1833 1012 1835 1015
rect 1843 1012 1845 1015
rect 1876 1012 1878 1015
rect 1919 1012 1921 1015
rect 1929 1012 1931 1015
rect 1962 1012 1964 1015
rect 2009 1012 2011 1015
rect 2019 1012 2021 1015
rect 2052 1012 2054 1015
rect 2104 1012 2106 1015
rect 2114 1012 2116 1015
rect 2147 1012 2149 1015
<< polycontact >>
rect 1612 3373 1616 3377
rect 1638 3373 1642 3377
rect 1664 3373 1668 3377
rect 1684 3373 1688 3377
rect 1774 3382 1778 3386
rect 1800 3382 1804 3386
rect 1826 3382 1830 3386
rect 1846 3382 1850 3386
rect 2011 3392 2015 3396
rect 1684 3358 1688 3362
rect 2037 3392 2041 3396
rect 2063 3392 2067 3396
rect 2083 3392 2087 3396
rect 1846 3367 1850 3371
rect 2083 3377 2087 3381
rect 1900 3277 1904 3281
rect 1910 3268 1914 3272
rect 1943 3277 1947 3281
rect 2028 3278 2032 3282
rect 2038 3269 2042 3273
rect 2071 3278 2075 3282
rect 2069 3205 2073 3209
rect 2079 3198 2083 3202
rect 2097 3200 2101 3204
rect 1621 3041 1625 3045
rect 1647 3041 1651 3045
rect 1673 3041 1677 3045
rect 1693 3041 1697 3045
rect 1783 3050 1787 3054
rect 1809 3050 1813 3054
rect 1835 3050 1839 3054
rect 1855 3050 1859 3054
rect 2020 3060 2024 3064
rect 1693 3026 1697 3030
rect 2046 3060 2050 3064
rect 2072 3060 2076 3064
rect 2092 3060 2096 3064
rect 1855 3035 1859 3039
rect 2092 3045 2096 3049
rect 1909 2945 1913 2949
rect 1919 2936 1923 2940
rect 1952 2945 1956 2949
rect 2037 2946 2041 2950
rect 2047 2937 2051 2941
rect 2080 2946 2084 2950
rect 2078 2873 2082 2877
rect 2088 2866 2092 2870
rect 2106 2868 2110 2872
rect 1642 2675 1646 2679
rect 1668 2675 1672 2679
rect 1694 2675 1698 2679
rect 1714 2675 1718 2679
rect 1804 2684 1808 2688
rect 1830 2684 1834 2688
rect 1856 2684 1860 2688
rect 1876 2684 1880 2688
rect 2041 2694 2045 2698
rect 1714 2660 1718 2664
rect 2067 2694 2071 2698
rect 2093 2694 2097 2698
rect 2113 2694 2117 2698
rect 1876 2669 1880 2673
rect 2113 2679 2117 2683
rect 1930 2579 1934 2583
rect 1940 2570 1944 2574
rect 1973 2579 1977 2583
rect 2058 2580 2062 2584
rect 2068 2571 2072 2575
rect 2101 2580 2105 2584
rect 2099 2507 2103 2511
rect 2109 2500 2113 2504
rect 2127 2502 2131 2506
rect 1670 2301 1674 2305
rect 1696 2301 1700 2305
rect 1722 2301 1726 2305
rect 1742 2301 1746 2305
rect 1832 2310 1836 2314
rect 1858 2310 1862 2314
rect 1884 2310 1888 2314
rect 1904 2310 1908 2314
rect 2069 2320 2073 2324
rect 1742 2286 1746 2290
rect 2095 2320 2099 2324
rect 2121 2320 2125 2324
rect 2141 2320 2145 2324
rect 1904 2295 1908 2299
rect 2141 2305 2145 2309
rect 1958 2205 1962 2209
rect 1968 2196 1972 2200
rect 2001 2205 2005 2209
rect 2086 2206 2090 2210
rect 2096 2197 2100 2201
rect 2129 2206 2133 2210
rect 2127 2133 2131 2137
rect 2137 2126 2141 2130
rect 2155 2128 2159 2132
rect 3955 1769 3959 1773
rect 3965 1762 3969 1766
rect 3975 1755 3979 1759
rect 3985 1748 3989 1752
rect 4016 1769 4020 1773
rect 1045 1711 1049 1715
rect 1101 1711 1105 1715
rect 1745 1695 1749 1699
rect 1755 1686 1759 1690
rect 1788 1695 1792 1699
rect 1831 1695 1835 1699
rect 1841 1686 1845 1690
rect 1874 1695 1878 1699
rect 1921 1695 1925 1699
rect 1931 1686 1935 1690
rect 1964 1695 1968 1699
rect 2016 1695 2020 1699
rect 2026 1686 2030 1690
rect 2059 1695 2063 1699
rect 2100 1695 2104 1699
rect 2110 1686 2114 1690
rect 2143 1695 2147 1699
rect 2186 1695 2190 1699
rect 2196 1686 2200 1690
rect 2229 1695 2233 1699
rect 2276 1695 2280 1699
rect 2286 1686 2290 1690
rect 2319 1695 2323 1699
rect 2371 1695 2375 1699
rect 2381 1686 2385 1690
rect 2414 1695 2418 1699
rect 1012 1634 1016 1638
rect 1022 1625 1026 1629
rect 1055 1634 1059 1638
rect 2960 1632 2964 1636
rect 2986 1632 2990 1636
rect 3012 1632 3016 1636
rect 3032 1632 3036 1636
rect 3096 1640 3100 1644
rect 3209 1632 3213 1636
rect 3032 1617 3036 1621
rect 3235 1632 3239 1636
rect 3261 1632 3265 1636
rect 3281 1632 3285 1636
rect 3345 1640 3349 1644
rect 3466 1632 3470 1636
rect 3281 1617 3285 1621
rect 3492 1632 3496 1636
rect 3518 1632 3522 1636
rect 3538 1632 3542 1636
rect 3602 1640 3606 1644
rect 3688 1632 3692 1636
rect 3538 1617 3542 1621
rect 3714 1632 3718 1636
rect 3740 1632 3744 1636
rect 3760 1632 3764 1636
rect 3824 1640 3828 1644
rect 3760 1617 3764 1621
rect 4254 1613 4258 1617
rect 4264 1606 4268 1610
rect 1318 1562 1322 1566
rect 1013 1549 1017 1553
rect 1023 1540 1027 1544
rect 1056 1549 1060 1553
rect 1328 1555 1332 1559
rect 1346 1557 1350 1561
rect 1013 1460 1017 1464
rect 1023 1451 1027 1455
rect 1056 1460 1060 1464
rect 1723 1451 1727 1455
rect 1733 1442 1737 1446
rect 1766 1451 1770 1455
rect 1809 1451 1813 1455
rect 1819 1442 1823 1446
rect 1852 1451 1856 1455
rect 1899 1451 1903 1455
rect 1909 1442 1913 1446
rect 1942 1451 1946 1455
rect 1994 1451 1998 1455
rect 2004 1442 2008 1446
rect 2037 1451 2041 1455
rect 2078 1451 2082 1455
rect 2088 1442 2092 1446
rect 2121 1451 2125 1455
rect 2164 1451 2168 1455
rect 2174 1442 2178 1446
rect 2207 1451 2211 1455
rect 2254 1451 2258 1455
rect 2264 1442 2268 1446
rect 2297 1451 2301 1455
rect 2349 1451 2353 1455
rect 2359 1442 2363 1446
rect 2392 1451 2396 1455
rect 3025 1443 3029 1447
rect 3035 1434 3039 1438
rect 3068 1443 3072 1447
rect 3227 1448 3231 1452
rect 3237 1441 3241 1445
rect 3247 1434 3251 1438
rect 3280 1448 3284 1452
rect 3482 1457 3486 1461
rect 3492 1450 3496 1454
rect 3502 1443 3506 1447
rect 3512 1436 3516 1440
rect 3543 1457 3547 1461
rect 3743 1467 3747 1471
rect 3753 1460 3757 1464
rect 3763 1453 3767 1457
rect 3773 1446 3777 1450
rect 3783 1438 3787 1442
rect 3816 1467 3820 1471
rect 4004 1395 4008 1399
rect 1013 1377 1017 1381
rect 1023 1368 1027 1372
rect 1056 1377 1060 1381
rect 4014 1388 4018 1392
rect 4024 1381 4028 1385
rect 4033 1374 4037 1378
rect 4052 1390 4056 1394
rect 3081 1282 3085 1286
rect 3137 1282 3141 1286
rect 3334 1282 3338 1286
rect 3597 1282 3601 1286
rect 1767 1134 1771 1138
rect 1777 1125 1781 1129
rect 1810 1134 1814 1138
rect 1853 1134 1857 1138
rect 1863 1125 1867 1129
rect 1896 1134 1900 1138
rect 1943 1134 1947 1138
rect 1953 1125 1957 1129
rect 1986 1134 1990 1138
rect 2038 1134 2042 1138
rect 2048 1125 2052 1129
rect 2081 1134 2085 1138
rect 2122 1134 2126 1138
rect 2132 1125 2136 1129
rect 2165 1134 2169 1138
rect 2208 1134 2212 1138
rect 2218 1125 2222 1129
rect 2251 1134 2255 1138
rect 2298 1134 2302 1138
rect 2308 1125 2312 1129
rect 2341 1134 2345 1138
rect 2393 1134 2397 1138
rect 2403 1125 2407 1129
rect 2436 1134 2440 1138
rect 1829 1033 1833 1037
rect 1839 1024 1843 1028
rect 1872 1033 1876 1037
rect 1915 1033 1919 1037
rect 1925 1024 1929 1028
rect 1958 1033 1962 1037
rect 2005 1033 2009 1037
rect 2015 1024 2019 1028
rect 2048 1033 2052 1037
rect 2100 1033 2104 1037
rect 2110 1024 2114 1028
rect 2143 1033 2147 1037
<< metal1 >>
rect 2293 3470 2301 3471
rect 2122 3464 2303 3470
rect 2122 3438 2127 3464
rect 1975 3434 2135 3438
rect 1975 3429 1980 3434
rect 1853 3428 1980 3429
rect 1739 3424 1980 3428
rect 1739 3419 1743 3424
rect 1605 3415 1743 3419
rect 1611 3402 1615 3415
rect 1627 3402 1631 3415
rect 1665 3402 1669 3415
rect 1685 3402 1689 3415
rect 1773 3411 1777 3424
rect 1789 3411 1793 3424
rect 1827 3411 1831 3424
rect 1847 3411 1851 3424
rect 2010 3421 2014 3434
rect 2026 3421 2030 3434
rect 2064 3421 2068 3434
rect 2084 3421 2088 3434
rect 1619 3377 1623 3396
rect 1646 3386 1650 3396
rect 1531 3373 1612 3377
rect 1619 3373 1638 3377
rect 1531 3364 1537 3373
rect 1586 3365 1605 3369
rect 1531 3282 1537 3359
rect 1619 3354 1623 3373
rect 1646 3354 1650 3381
rect 1677 3377 1681 3396
rect 1781 3386 1785 3405
rect 1808 3395 1812 3405
rect 1719 3385 1774 3386
rect 1712 3382 1774 3385
rect 1781 3382 1800 3386
rect 1712 3381 1748 3382
rect 1668 3373 1681 3377
rect 1677 3354 1681 3373
rect 1688 3370 1692 3377
rect 1719 3372 1725 3378
rect 1688 3358 1692 3365
rect 1611 3336 1615 3350
rect 1627 3336 1631 3350
rect 1665 3336 1669 3350
rect 1685 3336 1689 3350
rect 1606 3332 1691 3336
rect 1719 3282 1724 3336
rect 1530 3277 1725 3282
rect 1742 3281 1748 3381
rect 1760 3374 1767 3378
rect 1760 3373 1764 3374
rect 1781 3363 1785 3382
rect 1808 3363 1812 3390
rect 1839 3386 1843 3405
rect 1879 3394 1987 3396
rect 1874 3392 1987 3394
rect 2018 3396 2022 3415
rect 2045 3405 2049 3415
rect 1992 3392 2011 3396
rect 2018 3392 2037 3396
rect 1874 3390 1883 3392
rect 1830 3382 1843 3386
rect 1839 3363 1843 3382
rect 1850 3379 1854 3386
rect 1850 3367 1854 3374
rect 1980 3384 2004 3388
rect 1773 3345 1777 3359
rect 1789 3345 1793 3359
rect 1827 3345 1831 3359
rect 1847 3345 1851 3359
rect 1859 3345 1864 3347
rect 1768 3341 1864 3345
rect 1980 3335 1984 3384
rect 2018 3373 2022 3392
rect 2045 3373 2049 3400
rect 2076 3396 2080 3415
rect 2157 3400 2163 3405
rect 2067 3392 2080 3396
rect 2076 3373 2080 3392
rect 2087 3389 2091 3396
rect 2087 3377 2091 3384
rect 2010 3355 2014 3369
rect 2026 3355 2030 3369
rect 2064 3355 2068 3369
rect 2084 3355 2088 3369
rect 2010 3351 2254 3355
rect 1773 3331 1984 3335
rect 1893 3310 1957 3313
rect 1899 3295 1903 3310
rect 1918 3295 1922 3310
rect 1942 3295 1946 3310
rect 1908 3281 1912 3289
rect 1950 3281 1954 3289
rect 1980 3282 1984 3331
rect 2024 3311 2112 3314
rect 2027 3296 2031 3311
rect 2046 3296 2050 3311
rect 2070 3296 2074 3311
rect 2120 3311 2135 3314
rect 2036 3282 2040 3290
rect 2078 3282 2082 3290
rect 1960 3281 1973 3282
rect 1742 3277 1900 3281
rect 1908 3277 1943 3281
rect 1950 3277 1973 3281
rect 1980 3278 2028 3282
rect 2036 3278 2071 3282
rect 2078 3278 2135 3282
rect 1531 3045 1537 3277
rect 1743 3276 1892 3277
rect 1872 3268 1910 3272
rect 1918 3263 1922 3277
rect 1950 3263 1954 3277
rect 1869 3252 1894 3253
rect 1899 3252 1903 3259
rect 1942 3252 1946 3259
rect 1869 3249 1956 3252
rect 1966 3202 1973 3277
rect 1992 3269 2038 3273
rect 2046 3264 2050 3278
rect 2078 3264 2082 3278
rect 2027 3253 2031 3260
rect 2070 3253 2074 3260
rect 2024 3250 2089 3253
rect 2062 3236 2112 3241
rect 2068 3224 2072 3236
rect 2096 3224 2100 3236
rect 2022 3205 2069 3209
rect 2022 3161 2026 3205
rect 2086 3204 2090 3218
rect 2104 3204 2108 3218
rect 2065 3198 2079 3202
rect 2086 3200 2097 3204
rect 2104 3200 2120 3204
rect 2086 3194 2090 3200
rect 2077 3190 2090 3194
rect 2077 3186 2081 3190
rect 2104 3186 2108 3200
rect 2068 3175 2072 3182
rect 2086 3175 2090 3182
rect 2096 3175 2100 3182
rect 2064 3170 2113 3175
rect 2131 3161 2135 3278
rect 2022 3156 2135 3161
rect 2159 3147 2164 3205
rect 2248 3175 2254 3351
rect 1984 3102 2129 3106
rect 2134 3102 2144 3106
rect 1984 3097 1989 3102
rect 1862 3096 1989 3097
rect 1754 3092 1989 3096
rect 1754 3087 1758 3092
rect 1614 3083 1758 3087
rect 1620 3070 1624 3083
rect 1636 3070 1640 3083
rect 1674 3070 1678 3083
rect 1694 3070 1698 3083
rect 1782 3079 1786 3092
rect 1798 3079 1802 3092
rect 1836 3079 1840 3092
rect 1856 3079 1860 3092
rect 2019 3089 2023 3102
rect 2035 3089 2039 3102
rect 2073 3089 2077 3102
rect 2093 3089 2097 3102
rect 1628 3045 1632 3064
rect 1655 3054 1659 3064
rect 1531 3041 1621 3045
rect 1628 3041 1647 3045
rect 1531 2679 1537 3041
rect 1606 3033 1614 3037
rect 1628 3022 1632 3041
rect 1655 3022 1659 3049
rect 1686 3045 1690 3064
rect 1790 3054 1794 3073
rect 1817 3063 1821 3073
rect 1728 3053 1783 3054
rect 1721 3050 1783 3053
rect 1790 3050 1809 3054
rect 1721 3049 1757 3050
rect 1677 3041 1690 3045
rect 1686 3022 1690 3041
rect 1697 3038 1701 3045
rect 1728 3040 1734 3046
rect 1697 3026 1701 3033
rect 1620 3004 1624 3018
rect 1636 3004 1640 3018
rect 1674 3004 1678 3018
rect 1694 3004 1698 3018
rect 1615 3000 1703 3004
rect 1728 2998 1733 3004
rect 1751 2949 1757 3049
rect 1769 3042 1776 3046
rect 1769 3041 1773 3042
rect 1790 3031 1794 3050
rect 1817 3031 1821 3058
rect 1848 3054 1852 3073
rect 1888 3062 1996 3064
rect 1883 3060 1996 3062
rect 2027 3064 2031 3083
rect 2054 3073 2058 3083
rect 2001 3060 2020 3064
rect 2027 3060 2046 3064
rect 1883 3058 1892 3060
rect 1839 3050 1852 3054
rect 1848 3031 1852 3050
rect 1859 3047 1863 3054
rect 1859 3035 1863 3042
rect 1989 3052 2013 3056
rect 1782 3013 1786 3027
rect 1798 3013 1802 3027
rect 1836 3013 1840 3027
rect 1856 3013 1860 3027
rect 1868 3013 1873 3015
rect 1777 3009 1873 3013
rect 1989 3003 1993 3052
rect 2027 3041 2031 3060
rect 2054 3041 2058 3068
rect 2085 3064 2089 3083
rect 2166 3068 2172 3073
rect 2076 3060 2089 3064
rect 2085 3041 2089 3060
rect 2096 3057 2100 3064
rect 2096 3045 2100 3052
rect 2019 3023 2023 3037
rect 2035 3023 2039 3037
rect 2073 3023 2077 3037
rect 2093 3023 2097 3037
rect 2019 3019 2104 3023
rect 1782 2999 1993 3003
rect 1902 2978 1966 2981
rect 1908 2963 1912 2978
rect 1927 2963 1931 2978
rect 1951 2963 1955 2978
rect 1917 2949 1921 2957
rect 1959 2949 1963 2957
rect 1989 2950 1993 2999
rect 2033 2979 2121 2982
rect 2036 2964 2040 2979
rect 2055 2964 2059 2979
rect 2079 2964 2083 2979
rect 2129 2979 2144 2982
rect 2045 2950 2049 2958
rect 2087 2950 2091 2958
rect 1969 2949 1982 2950
rect 1751 2945 1909 2949
rect 1917 2945 1952 2949
rect 1959 2945 1982 2949
rect 1989 2946 2037 2950
rect 2045 2946 2080 2950
rect 2087 2946 2144 2950
rect 1752 2944 1910 2945
rect 1881 2936 1919 2940
rect 1927 2931 1931 2945
rect 1959 2931 1963 2945
rect 1878 2920 1903 2921
rect 1908 2920 1912 2927
rect 1951 2920 1955 2927
rect 1878 2917 1965 2920
rect 1975 2870 1982 2945
rect 2001 2937 2047 2941
rect 2055 2932 2059 2946
rect 2087 2932 2091 2946
rect 2036 2921 2040 2928
rect 2079 2921 2083 2928
rect 2033 2918 2098 2921
rect 2071 2904 2121 2909
rect 2077 2892 2081 2904
rect 2105 2892 2109 2904
rect 2031 2873 2078 2877
rect 2031 2829 2035 2873
rect 2095 2872 2099 2886
rect 2113 2872 2117 2886
rect 2074 2866 2088 2870
rect 2095 2868 2106 2872
rect 2113 2868 2129 2872
rect 2095 2862 2099 2868
rect 2086 2858 2099 2862
rect 2086 2854 2090 2858
rect 2113 2854 2117 2868
rect 2077 2843 2081 2850
rect 2095 2843 2099 2850
rect 2105 2843 2109 2850
rect 2073 2838 2127 2843
rect 2140 2829 2144 2946
rect 2031 2824 2144 2829
rect 2168 2781 2173 2873
rect 2248 2843 2254 3170
rect 2293 3121 2301 3464
rect 2145 2740 2149 2745
rect 2005 2736 2165 2740
rect 2005 2731 2010 2736
rect 1883 2730 2010 2731
rect 1777 2726 2010 2730
rect 1778 2721 1782 2726
rect 1635 2717 1782 2721
rect 1641 2704 1645 2717
rect 1657 2704 1661 2717
rect 1695 2704 1699 2717
rect 1715 2704 1719 2717
rect 1803 2713 1807 2726
rect 1819 2713 1823 2726
rect 1857 2713 1861 2726
rect 1877 2713 1881 2726
rect 2040 2723 2044 2736
rect 2056 2723 2060 2736
rect 2094 2723 2098 2736
rect 2114 2723 2118 2736
rect 1649 2679 1653 2698
rect 1676 2688 1680 2698
rect 1530 2675 1642 2679
rect 1649 2675 1668 2679
rect 1211 1790 1217 2525
rect 1531 2297 1537 2675
rect 1631 2667 1635 2671
rect 1649 2656 1653 2675
rect 1676 2656 1680 2683
rect 1707 2679 1711 2698
rect 1811 2688 1815 2707
rect 1838 2697 1842 2707
rect 1749 2687 1804 2688
rect 1742 2684 1804 2687
rect 1811 2684 1830 2688
rect 1742 2683 1778 2684
rect 1698 2675 1711 2679
rect 1707 2656 1711 2675
rect 1718 2672 1722 2679
rect 1718 2660 1722 2667
rect 1737 2674 1755 2680
rect 1641 2638 1645 2652
rect 1657 2638 1661 2652
rect 1695 2638 1699 2652
rect 1715 2638 1719 2652
rect 1636 2634 1722 2638
rect 1737 2530 1743 2674
rect 1749 2632 1754 2638
rect 1772 2583 1778 2683
rect 1790 2676 1797 2680
rect 1790 2675 1794 2676
rect 1811 2665 1815 2684
rect 1838 2665 1842 2692
rect 1869 2688 1873 2707
rect 1909 2696 2017 2698
rect 1904 2694 2017 2696
rect 2048 2698 2052 2717
rect 2075 2707 2079 2717
rect 2022 2694 2041 2698
rect 2048 2694 2067 2698
rect 1904 2692 1913 2694
rect 1860 2684 1873 2688
rect 1869 2665 1873 2684
rect 1880 2681 1884 2688
rect 1880 2669 1884 2676
rect 2010 2686 2034 2690
rect 1803 2647 1807 2661
rect 1819 2647 1823 2661
rect 1857 2647 1861 2661
rect 1877 2647 1881 2661
rect 1889 2647 1894 2649
rect 1798 2643 1894 2647
rect 2010 2637 2014 2686
rect 2048 2675 2052 2694
rect 2075 2675 2079 2702
rect 2106 2698 2110 2717
rect 2187 2702 2193 2707
rect 2097 2694 2110 2698
rect 2106 2675 2110 2694
rect 2117 2691 2121 2698
rect 2117 2679 2121 2686
rect 2040 2657 2044 2671
rect 2056 2657 2060 2671
rect 2094 2657 2098 2671
rect 2114 2657 2118 2671
rect 2040 2653 2125 2657
rect 1803 2633 2014 2637
rect 1923 2612 1987 2615
rect 1929 2597 1933 2612
rect 1948 2597 1952 2612
rect 1972 2597 1976 2612
rect 1938 2583 1942 2591
rect 1980 2583 1984 2591
rect 2010 2584 2014 2633
rect 2054 2613 2142 2616
rect 2057 2598 2061 2613
rect 2076 2598 2080 2613
rect 2100 2598 2104 2613
rect 2150 2613 2165 2616
rect 2066 2584 2070 2592
rect 2108 2584 2112 2592
rect 1990 2583 2003 2584
rect 1772 2579 1930 2583
rect 1938 2579 1973 2583
rect 1980 2579 2003 2583
rect 2010 2580 2058 2584
rect 2066 2580 2101 2584
rect 2108 2580 2165 2584
rect 1773 2578 1922 2579
rect 1902 2570 1940 2574
rect 1948 2565 1952 2579
rect 1980 2565 1984 2579
rect 1899 2554 1924 2555
rect 1929 2554 1933 2561
rect 1972 2554 1976 2561
rect 1899 2551 1986 2554
rect 1996 2504 2003 2579
rect 2022 2571 2068 2575
rect 2076 2566 2080 2580
rect 2108 2566 2112 2580
rect 2057 2555 2061 2562
rect 2100 2555 2104 2562
rect 2054 2552 2119 2555
rect 2092 2538 2142 2543
rect 2098 2526 2102 2538
rect 2126 2526 2130 2538
rect 2052 2507 2099 2511
rect 2052 2463 2056 2507
rect 2116 2506 2120 2520
rect 2134 2506 2138 2520
rect 2095 2500 2109 2504
rect 2116 2502 2127 2506
rect 2134 2502 2150 2506
rect 2116 2496 2120 2502
rect 2107 2492 2120 2496
rect 2107 2488 2111 2492
rect 2134 2488 2138 2502
rect 2098 2477 2102 2484
rect 2116 2477 2120 2484
rect 2126 2477 2130 2484
rect 2094 2472 2148 2477
rect 2161 2463 2165 2580
rect 2052 2458 2165 2463
rect 2189 2411 2194 2507
rect 2248 2478 2254 2838
rect 2033 2362 2173 2366
rect 2178 2362 2193 2366
rect 2033 2357 2038 2362
rect 1911 2356 2038 2357
rect 1788 2352 2038 2356
rect 1788 2347 1793 2352
rect 1663 2343 1793 2347
rect 1669 2330 1673 2343
rect 1685 2330 1689 2343
rect 1723 2330 1727 2343
rect 1743 2330 1747 2343
rect 1831 2339 1835 2352
rect 1847 2339 1851 2352
rect 1885 2339 1889 2352
rect 1905 2339 1909 2352
rect 2068 2349 2072 2362
rect 2084 2349 2088 2362
rect 2122 2349 2126 2362
rect 2142 2349 2146 2362
rect 1607 2307 1659 2310
rect 1655 2305 1659 2307
rect 1677 2305 1681 2324
rect 1704 2314 1708 2324
rect 1655 2301 1670 2305
rect 1677 2301 1696 2305
rect 1267 2293 1663 2297
rect 1267 2292 1537 2293
rect 1531 2291 1537 2292
rect 1677 2282 1681 2301
rect 1704 2282 1708 2309
rect 1735 2305 1739 2324
rect 1839 2314 1843 2333
rect 1866 2323 1870 2333
rect 1777 2313 1832 2314
rect 1770 2310 1832 2313
rect 1839 2310 1858 2314
rect 1770 2309 1806 2310
rect 1726 2301 1739 2305
rect 1735 2282 1739 2301
rect 1746 2298 1750 2305
rect 1746 2286 1750 2293
rect 1766 2300 1783 2306
rect 1669 2264 1673 2278
rect 1685 2264 1689 2278
rect 1723 2264 1727 2278
rect 1743 2264 1747 2278
rect 1664 2260 1750 2264
rect 1766 2164 1771 2300
rect 1777 2258 1782 2264
rect 1800 2209 1806 2309
rect 1818 2302 1825 2306
rect 1818 2301 1822 2302
rect 1839 2291 1843 2310
rect 1866 2291 1870 2318
rect 1897 2314 1901 2333
rect 1937 2322 2045 2324
rect 1932 2320 2045 2322
rect 2076 2324 2080 2343
rect 2103 2333 2107 2343
rect 2050 2320 2069 2324
rect 2076 2320 2095 2324
rect 1932 2318 1941 2320
rect 1888 2310 1901 2314
rect 1897 2291 1901 2310
rect 1908 2307 1912 2314
rect 1908 2295 1912 2302
rect 2038 2312 2062 2316
rect 1831 2273 1835 2287
rect 1847 2273 1851 2287
rect 1885 2273 1889 2287
rect 1905 2273 1909 2287
rect 1917 2273 1922 2275
rect 1826 2269 1922 2273
rect 2038 2263 2042 2312
rect 2076 2301 2080 2320
rect 2103 2301 2107 2328
rect 2134 2324 2138 2343
rect 2215 2328 2221 2333
rect 2125 2320 2138 2324
rect 2134 2301 2138 2320
rect 2145 2317 2149 2324
rect 2145 2305 2149 2312
rect 2068 2283 2072 2297
rect 2084 2283 2088 2297
rect 2122 2283 2126 2297
rect 2142 2283 2146 2297
rect 2068 2279 2153 2283
rect 1831 2259 2042 2263
rect 1951 2238 2015 2241
rect 1957 2223 1961 2238
rect 1976 2223 1980 2238
rect 2000 2223 2004 2238
rect 1966 2209 1970 2217
rect 2008 2209 2012 2217
rect 2038 2210 2042 2259
rect 2082 2239 2170 2242
rect 2085 2224 2089 2239
rect 2104 2224 2108 2239
rect 2128 2224 2132 2239
rect 2178 2239 2193 2242
rect 2094 2210 2098 2218
rect 2136 2210 2140 2218
rect 2018 2209 2031 2210
rect 1800 2205 1958 2209
rect 1966 2205 2001 2209
rect 2008 2205 2031 2209
rect 2038 2206 2086 2210
rect 2094 2206 2129 2210
rect 2136 2206 2193 2210
rect 1801 2204 1950 2205
rect 1930 2196 1968 2200
rect 1976 2191 1980 2205
rect 2008 2191 2012 2205
rect 1928 2180 1952 2181
rect 1957 2180 1961 2187
rect 2000 2180 2004 2187
rect 1928 2177 2014 2180
rect 1766 2158 1804 2164
rect 1799 2099 1804 2158
rect 2024 2130 2031 2205
rect 2050 2197 2096 2201
rect 2104 2192 2108 2206
rect 2136 2192 2140 2206
rect 2085 2181 2089 2188
rect 2128 2181 2132 2188
rect 2082 2178 2147 2181
rect 2120 2164 2170 2169
rect 2126 2152 2130 2164
rect 2154 2152 2158 2164
rect 2080 2133 2127 2137
rect 2080 2089 2084 2133
rect 2144 2132 2148 2146
rect 2162 2132 2166 2146
rect 2123 2126 2137 2130
rect 2144 2128 2155 2132
rect 2162 2128 2178 2132
rect 2144 2122 2148 2128
rect 2135 2118 2148 2122
rect 2135 2114 2139 2118
rect 2162 2114 2166 2128
rect 2126 2103 2130 2110
rect 2144 2103 2148 2110
rect 2154 2103 2158 2110
rect 2122 2098 2168 2103
rect 2189 2089 2193 2206
rect 2217 2128 2222 2133
rect 2248 2103 2254 2472
rect 2293 2750 2301 3116
rect 2293 2384 2301 2745
rect 2609 2384 2615 2386
rect 2293 2383 2615 2384
rect 2301 2378 2615 2383
rect 2255 2098 2525 2103
rect 2248 2097 2532 2098
rect 2080 2084 2193 2089
rect 1569 1799 2073 1804
rect 2157 1792 2163 1908
rect 2250 1812 2471 1819
rect 1211 1785 1983 1790
rect 2340 1789 2379 1797
rect 1211 1784 1792 1785
rect 2609 1778 2615 2378
rect 2485 1774 2615 1778
rect 2486 1761 2491 1774
rect 1148 1739 1318 1742
rect 1148 1738 1153 1739
rect 1042 1733 1148 1736
rect 1049 1727 1052 1733
rect 1105 1727 1108 1733
rect 1148 1730 1153 1733
rect 955 1711 1045 1715
rect 1056 1714 1059 1723
rect 1056 1711 1063 1714
rect 955 1553 959 1711
rect 1056 1707 1059 1711
rect 1095 1711 1101 1715
rect 1112 1714 1115 1723
rect 1112 1711 1127 1714
rect 1112 1707 1115 1711
rect 1049 1699 1052 1703
rect 1105 1699 1108 1703
rect 1042 1696 1119 1699
rect 1005 1667 1148 1670
rect 1011 1652 1015 1667
rect 1030 1652 1034 1667
rect 1054 1652 1058 1667
rect 1020 1638 1024 1646
rect 1062 1638 1066 1646
rect 968 1634 1012 1638
rect 1020 1634 1055 1638
rect 1062 1634 1229 1638
rect 993 1625 1022 1629
rect 1030 1620 1034 1634
rect 1062 1620 1066 1634
rect 1011 1609 1015 1616
rect 1054 1609 1058 1616
rect 1004 1606 1119 1609
rect 1119 1585 1124 1586
rect 1006 1582 1148 1585
rect 1012 1567 1016 1582
rect 1031 1567 1035 1582
rect 1055 1567 1059 1582
rect 1119 1581 1124 1582
rect 1225 1566 1229 1634
rect 1313 1598 1318 1739
rect 1679 1739 1727 1744
rect 1311 1593 1368 1598
rect 1317 1581 1321 1593
rect 1345 1581 1349 1593
rect 1225 1562 1318 1566
rect 1021 1553 1025 1561
rect 1063 1553 1067 1561
rect 1335 1561 1339 1575
rect 1353 1561 1357 1575
rect 1679 1561 1683 1739
rect 2486 1731 2490 1761
rect 1738 1728 2490 1731
rect 1744 1713 1748 1728
rect 1763 1713 1767 1728
rect 1787 1713 1791 1728
rect 1830 1713 1834 1728
rect 1849 1713 1853 1728
rect 1873 1713 1877 1728
rect 1920 1713 1924 1728
rect 1939 1713 1943 1728
rect 1963 1713 1967 1728
rect 2015 1713 2019 1728
rect 2034 1713 2038 1728
rect 2058 1713 2062 1728
rect 2099 1713 2103 1728
rect 2118 1713 2122 1728
rect 2142 1713 2146 1728
rect 2185 1713 2189 1728
rect 2204 1713 2208 1728
rect 2228 1713 2232 1728
rect 2275 1713 2279 1728
rect 2294 1713 2298 1728
rect 2318 1713 2322 1728
rect 2370 1713 2374 1728
rect 2389 1713 2393 1728
rect 2413 1713 2417 1728
rect 1753 1699 1757 1707
rect 1710 1695 1745 1699
rect 1753 1695 1788 1699
rect 1733 1686 1755 1690
rect 1763 1681 1767 1695
rect 1795 1681 1799 1707
rect 1839 1699 1843 1707
rect 1881 1699 1885 1707
rect 1929 1699 1933 1707
rect 1971 1699 1975 1707
rect 2024 1699 2028 1707
rect 2066 1699 2070 1707
rect 2108 1699 2112 1707
rect 2150 1699 2154 1707
rect 2194 1699 2198 1707
rect 2236 1699 2240 1707
rect 2284 1699 2288 1707
rect 2326 1699 2330 1707
rect 2379 1699 2383 1707
rect 2421 1699 2425 1707
rect 1804 1695 1808 1699
rect 1819 1695 1823 1699
rect 1828 1695 1831 1699
rect 1839 1695 1874 1699
rect 1881 1695 1890 1699
rect 1818 1686 1841 1690
rect 1849 1681 1853 1695
rect 1881 1681 1885 1695
rect 1909 1695 1913 1699
rect 1918 1695 1921 1699
rect 1929 1695 1964 1699
rect 1971 1695 1983 1699
rect 1908 1686 1931 1690
rect 1939 1681 1943 1695
rect 1971 1681 1975 1695
rect 2004 1695 2008 1699
rect 2013 1695 2016 1699
rect 2024 1695 2059 1699
rect 2066 1695 2073 1699
rect 2002 1686 2026 1690
rect 2034 1681 2038 1695
rect 2066 1681 2070 1695
rect 2078 1695 2079 1699
rect 2088 1695 2092 1699
rect 2097 1695 2100 1699
rect 2108 1695 2143 1699
rect 2150 1695 2157 1699
rect 2088 1686 2110 1690
rect 2118 1681 2122 1695
rect 2150 1681 2154 1695
rect 2162 1695 2163 1699
rect 2174 1695 2178 1699
rect 2183 1695 2186 1699
rect 2194 1695 2229 1699
rect 2236 1695 2243 1699
rect 2173 1686 2196 1690
rect 2204 1681 2208 1695
rect 2236 1681 2240 1695
rect 2248 1695 2249 1699
rect 2264 1695 2268 1699
rect 2273 1695 2276 1699
rect 2284 1695 2319 1699
rect 2326 1695 2334 1699
rect 2263 1686 2286 1690
rect 2294 1681 2298 1695
rect 2326 1681 2330 1695
rect 2359 1695 2363 1699
rect 2368 1695 2371 1699
rect 2379 1695 2414 1699
rect 2421 1695 2429 1699
rect 2357 1686 2381 1690
rect 2389 1681 2393 1695
rect 2421 1681 2425 1695
rect 1744 1670 1748 1677
rect 1787 1670 1791 1677
rect 1830 1670 1834 1677
rect 1873 1670 1877 1677
rect 1920 1670 1924 1677
rect 1963 1670 1967 1677
rect 2015 1670 2019 1677
rect 2058 1670 2062 1677
rect 2099 1670 2103 1677
rect 2142 1670 2146 1677
rect 2185 1670 2189 1677
rect 2228 1670 2232 1677
rect 2275 1670 2279 1677
rect 2318 1670 2322 1677
rect 2370 1670 2374 1677
rect 2413 1670 2417 1677
rect 1737 1667 2429 1670
rect 1295 1555 1328 1559
rect 1335 1557 1346 1561
rect 1353 1557 1683 1561
rect 955 1549 1013 1553
rect 1021 1549 1056 1553
rect 1063 1549 1261 1553
rect 1295 1553 1299 1555
rect 1266 1549 1299 1553
rect 1335 1551 1339 1557
rect 955 1381 959 1549
rect 993 1540 1023 1544
rect 1031 1535 1035 1549
rect 1063 1535 1067 1549
rect 1326 1547 1339 1551
rect 1326 1543 1330 1547
rect 1353 1543 1357 1557
rect 1012 1524 1016 1531
rect 1055 1524 1059 1531
rect 1317 1532 1321 1539
rect 1335 1532 1339 1539
rect 1345 1532 1349 1539
rect 1139 1527 1367 1532
rect 1005 1521 1119 1524
rect 1006 1493 1148 1496
rect 1657 1495 1705 1500
rect 1012 1478 1016 1493
rect 1031 1478 1035 1493
rect 1055 1478 1059 1493
rect 1021 1464 1025 1472
rect 1063 1464 1067 1472
rect 1657 1464 1661 1495
rect 2486 1487 2490 1728
rect 1716 1484 2490 1487
rect 968 1460 1013 1464
rect 1021 1460 1056 1464
rect 1063 1460 1661 1464
rect 1722 1469 1726 1484
rect 1741 1469 1745 1484
rect 1765 1469 1769 1484
rect 1808 1469 1812 1484
rect 1827 1469 1831 1484
rect 1851 1469 1855 1484
rect 1898 1469 1902 1484
rect 1917 1469 1921 1484
rect 1941 1469 1945 1484
rect 1993 1469 1997 1484
rect 2012 1469 2016 1484
rect 2036 1469 2040 1484
rect 2077 1469 2081 1484
rect 2096 1469 2100 1484
rect 2120 1469 2124 1484
rect 2163 1469 2167 1484
rect 2182 1469 2186 1484
rect 2206 1469 2210 1484
rect 2253 1469 2257 1484
rect 2272 1469 2276 1484
rect 2296 1469 2300 1484
rect 2348 1469 2352 1484
rect 2367 1469 2371 1484
rect 2391 1469 2395 1484
rect 980 1451 1023 1455
rect 1031 1446 1035 1460
rect 1063 1446 1067 1460
rect 1731 1455 1735 1463
rect 1773 1455 1777 1463
rect 1817 1455 1821 1463
rect 1859 1455 1863 1463
rect 1907 1455 1911 1463
rect 1949 1455 1953 1463
rect 2002 1455 2006 1463
rect 2044 1455 2048 1463
rect 2086 1455 2090 1463
rect 2128 1455 2132 1463
rect 2172 1455 2176 1463
rect 2214 1455 2218 1463
rect 2262 1455 2266 1463
rect 2304 1455 2308 1463
rect 2357 1455 2361 1463
rect 2399 1455 2403 1463
rect 1686 1451 1723 1455
rect 1731 1451 1766 1455
rect 1773 1451 1781 1455
rect 1012 1435 1016 1442
rect 1055 1435 1059 1442
rect 1711 1442 1733 1446
rect 1741 1437 1745 1451
rect 1773 1437 1777 1451
rect 1797 1451 1801 1455
rect 1806 1451 1809 1455
rect 1817 1451 1852 1455
rect 1859 1451 1867 1455
rect 1796 1442 1819 1446
rect 1827 1437 1831 1451
rect 1859 1437 1863 1451
rect 1887 1451 1891 1455
rect 1896 1451 1899 1455
rect 1907 1451 1942 1455
rect 1949 1451 1958 1455
rect 1886 1442 1909 1446
rect 1917 1437 1921 1451
rect 1949 1437 1953 1451
rect 1982 1451 1986 1455
rect 1991 1451 1994 1455
rect 2002 1451 2037 1455
rect 2044 1451 2051 1455
rect 1980 1442 2004 1446
rect 2012 1437 2016 1451
rect 2044 1437 2048 1451
rect 2056 1451 2057 1455
rect 2066 1451 2070 1455
rect 2075 1451 2078 1455
rect 2086 1451 2121 1455
rect 2128 1451 2135 1455
rect 2066 1442 2088 1446
rect 2096 1437 2100 1451
rect 2128 1437 2132 1451
rect 2140 1451 2141 1455
rect 2152 1451 2156 1455
rect 2161 1451 2164 1455
rect 2172 1451 2207 1455
rect 2214 1451 2221 1455
rect 2151 1442 2174 1446
rect 2182 1437 2186 1451
rect 2214 1437 2218 1451
rect 2226 1451 2227 1455
rect 2242 1451 2246 1455
rect 2251 1451 2254 1455
rect 2262 1451 2297 1455
rect 2304 1451 2311 1455
rect 2241 1442 2264 1446
rect 2272 1437 2276 1451
rect 2304 1437 2308 1451
rect 2316 1451 2317 1455
rect 2337 1451 2341 1455
rect 2346 1451 2349 1455
rect 2357 1451 2392 1455
rect 2399 1451 2407 1455
rect 2335 1442 2359 1446
rect 2367 1437 2371 1451
rect 2399 1437 2403 1451
rect 1005 1432 1119 1435
rect 1722 1426 1726 1433
rect 1765 1426 1769 1433
rect 1808 1426 1812 1433
rect 1851 1426 1855 1433
rect 1898 1426 1902 1433
rect 1941 1426 1945 1433
rect 1993 1426 1997 1433
rect 2036 1426 2040 1433
rect 2077 1426 2081 1433
rect 2120 1426 2124 1433
rect 2163 1426 2167 1433
rect 2206 1426 2210 1433
rect 2253 1426 2257 1433
rect 2296 1426 2300 1433
rect 2348 1426 2352 1433
rect 2391 1426 2395 1433
rect 1715 1423 2405 1426
rect 1006 1410 1148 1413
rect 1012 1395 1016 1410
rect 1031 1395 1035 1410
rect 1055 1395 1059 1410
rect 1786 1408 2434 1412
rect 1021 1381 1025 1389
rect 1063 1381 1067 1389
rect 955 1377 1013 1381
rect 1021 1377 1056 1381
rect 1063 1377 1323 1381
rect 1872 1380 2434 1385
rect 980 1368 1023 1372
rect 1031 1363 1035 1377
rect 1063 1363 1067 1377
rect 1012 1352 1016 1359
rect 1055 1352 1059 1359
rect 1005 1349 1119 1352
rect 1315 1222 1323 1377
rect 1963 1356 2436 1361
rect 2056 1343 2436 1348
rect 2140 1320 2436 1325
rect 2226 1301 2438 1306
rect 2221 1300 2438 1301
rect 2316 1291 2454 1296
rect 1315 1183 1322 1222
rect 1315 1178 1749 1183
rect 2486 1171 2490 1484
rect 2641 1349 2650 1715
rect 2667 1326 2675 1811
rect 2736 1794 2744 1854
rect 3948 1805 4326 1806
rect 3948 1802 4448 1805
rect 2710 1307 2720 1742
rect 2737 1296 2744 1794
rect 2795 1456 2803 1788
rect 3954 1787 3958 1802
rect 3973 1787 3977 1802
rect 3993 1787 3997 1802
rect 4015 1787 4019 1802
rect 4320 1799 4448 1802
rect 3963 1773 3967 1781
rect 3983 1773 3987 1781
rect 4023 1773 4027 1781
rect 3151 1769 3955 1773
rect 3963 1769 4016 1773
rect 4023 1769 4139 1773
rect 3399 1762 3965 1766
rect 3644 1755 3975 1759
rect 3892 1748 3985 1752
rect 2872 1689 2940 1696
rect 2873 1385 2880 1689
rect 2953 1674 3820 1678
rect 2959 1661 2963 1674
rect 2975 1661 2979 1674
rect 3013 1661 3017 1674
rect 3033 1661 3037 1674
rect 3093 1665 3096 1674
rect 3093 1662 3118 1665
rect 3100 1656 3103 1662
rect 3208 1661 3212 1674
rect 3224 1661 3228 1674
rect 3262 1661 3266 1674
rect 3282 1661 3286 1674
rect 3342 1665 3345 1674
rect 3342 1662 3367 1665
rect 2967 1636 2971 1655
rect 2994 1645 2998 1655
rect 2917 1632 2960 1636
rect 2967 1632 2986 1636
rect 2917 1457 2923 1632
rect 2946 1624 2953 1628
rect 2946 1623 2950 1624
rect 2967 1613 2971 1632
rect 2994 1613 2998 1640
rect 3025 1636 3029 1655
rect 3349 1656 3352 1662
rect 3465 1661 3469 1674
rect 3481 1661 3485 1674
rect 3519 1661 3523 1674
rect 3539 1661 3543 1674
rect 3599 1665 3602 1674
rect 3599 1662 3624 1665
rect 3060 1640 3096 1644
rect 3107 1643 3110 1652
rect 3107 1640 3144 1643
rect 3107 1636 3110 1640
rect 3216 1636 3220 1655
rect 3243 1645 3247 1655
rect 3016 1632 3029 1636
rect 3025 1613 3029 1632
rect 3036 1629 3040 1636
rect 3100 1628 3103 1632
rect 3167 1632 3209 1636
rect 3216 1632 3235 1636
rect 3036 1617 3040 1624
rect 3093 1625 3123 1628
rect 2959 1595 2963 1609
rect 2975 1595 2979 1609
rect 3013 1595 3017 1609
rect 3033 1595 3037 1609
rect 3093 1595 3096 1625
rect 3177 1624 3202 1628
rect 3216 1613 3220 1632
rect 3243 1613 3247 1640
rect 3274 1636 3278 1655
rect 3606 1656 3609 1662
rect 3687 1661 3691 1674
rect 3703 1661 3707 1674
rect 3741 1661 3745 1674
rect 3761 1661 3765 1674
rect 3821 1665 3824 1674
rect 3821 1662 3846 1665
rect 3309 1640 3345 1644
rect 3356 1643 3359 1652
rect 3356 1640 3393 1643
rect 3356 1636 3359 1640
rect 3473 1636 3477 1655
rect 3500 1645 3504 1655
rect 3265 1632 3278 1636
rect 3274 1613 3278 1632
rect 3285 1629 3289 1636
rect 3349 1628 3352 1632
rect 3443 1632 3466 1636
rect 3473 1632 3492 1636
rect 3285 1617 3289 1624
rect 3342 1625 3367 1628
rect 3208 1595 3212 1609
rect 3224 1595 3228 1609
rect 3262 1595 3266 1609
rect 3282 1595 3286 1609
rect 3342 1595 3345 1625
rect 3419 1624 3459 1628
rect 3473 1613 3477 1632
rect 3500 1613 3504 1640
rect 3531 1636 3535 1655
rect 3828 1656 3831 1662
rect 3566 1640 3602 1644
rect 3613 1643 3616 1652
rect 3613 1640 3637 1643
rect 3613 1636 3616 1640
rect 3695 1636 3699 1655
rect 3722 1645 3726 1655
rect 3522 1632 3535 1636
rect 3531 1613 3535 1632
rect 3542 1629 3546 1636
rect 3606 1628 3609 1632
rect 3663 1632 3688 1636
rect 3695 1632 3714 1636
rect 3542 1617 3546 1624
rect 3599 1625 3624 1628
rect 3465 1595 3469 1609
rect 3481 1595 3485 1609
rect 3519 1595 3523 1609
rect 3539 1595 3543 1609
rect 3599 1595 3602 1625
rect 3677 1624 3681 1628
rect 3695 1613 3699 1632
rect 3722 1613 3726 1640
rect 3753 1636 3757 1655
rect 3788 1640 3824 1644
rect 3835 1643 3838 1652
rect 3892 1643 3896 1748
rect 3993 1744 3997 1769
rect 4023 1744 4027 1769
rect 3954 1733 3958 1740
rect 4015 1733 4019 1740
rect 3947 1730 4028 1733
rect 3835 1640 3896 1643
rect 3835 1636 3838 1640
rect 3744 1632 3757 1636
rect 3753 1613 3757 1632
rect 3764 1629 3768 1636
rect 3828 1628 3831 1632
rect 3764 1617 3768 1624
rect 3821 1625 3847 1628
rect 3687 1595 3691 1609
rect 3703 1595 3707 1609
rect 3741 1595 3745 1609
rect 3761 1595 3765 1609
rect 3821 1595 3824 1625
rect 2954 1592 3824 1595
rect 3843 1552 3847 1625
rect 4134 1617 4139 1769
rect 4320 1681 4326 1799
rect 4320 1649 4326 1674
rect 4247 1644 4326 1649
rect 4253 1632 4257 1644
rect 4134 1613 4254 1617
rect 4271 1612 4275 1626
rect 4134 1606 4264 1610
rect 4271 1608 4283 1612
rect 3316 1524 3598 1529
rect 3647 1500 3826 1504
rect 3647 1493 3651 1500
rect 3370 1490 3651 1493
rect 3371 1485 3376 1490
rect 3190 1481 3376 1485
rect 3190 1479 3194 1481
rect 3018 1476 3194 1479
rect 3024 1461 3028 1476
rect 3043 1461 3047 1476
rect 2917 1453 3013 1457
rect 3067 1461 3071 1476
rect 3226 1466 3230 1481
rect 3245 1466 3249 1481
rect 3279 1466 3283 1481
rect 3481 1475 3485 1490
rect 3500 1475 3504 1490
rect 3520 1475 3524 1490
rect 3542 1475 3546 1490
rect 3742 1485 3746 1500
rect 3761 1485 3765 1500
rect 3781 1485 3785 1500
rect 3815 1485 3819 1500
rect 3150 1462 3209 1465
rect 2917 1414 2925 1453
rect 3009 1447 3013 1453
rect 3033 1447 3037 1455
rect 3075 1447 3079 1455
rect 3205 1452 3209 1462
rect 3235 1452 3239 1460
rect 3255 1452 3259 1460
rect 3287 1452 3291 1460
rect 3490 1461 3494 1469
rect 3510 1461 3514 1469
rect 3550 1461 3554 1469
rect 3751 1471 3755 1479
rect 3771 1471 3775 1479
rect 3791 1471 3795 1479
rect 3823 1471 3827 1479
rect 3604 1467 3743 1471
rect 3751 1467 3816 1471
rect 3823 1467 3874 1471
rect 3423 1457 3482 1461
rect 3490 1457 3543 1461
rect 3550 1457 3576 1461
rect 3205 1448 3227 1452
rect 3235 1448 3280 1452
rect 3287 1448 3344 1452
rect 3009 1443 3025 1447
rect 3033 1443 3068 1447
rect 3075 1443 3095 1447
rect 2992 1434 3035 1438
rect 3043 1429 3047 1443
rect 3075 1429 3079 1443
rect 3172 1441 3237 1445
rect 3185 1436 3247 1438
rect 3190 1434 3247 1436
rect 3255 1431 3259 1448
rect 3287 1431 3291 1448
rect 3440 1450 3492 1454
rect 3447 1443 3502 1447
rect 3447 1438 3451 1443
rect 3375 1435 3451 1438
rect 3470 1436 3512 1440
rect 3470 1431 3474 1436
rect 3520 1432 3524 1457
rect 3550 1432 3554 1457
rect 3633 1460 3753 1464
rect 3650 1453 3763 1457
rect 3665 1446 3773 1450
rect 3665 1445 3728 1446
rect 3731 1438 3783 1442
rect 3731 1436 3736 1438
rect 3024 1418 3028 1425
rect 3067 1418 3071 1425
rect 3226 1420 3230 1427
rect 3279 1420 3283 1427
rect 3444 1427 3474 1431
rect 3791 1435 3795 1467
rect 3823 1435 3827 1467
rect 3481 1421 3485 1428
rect 3542 1421 3546 1428
rect 3742 1424 3746 1431
rect 3815 1424 3819 1431
rect 4069 1430 4074 1500
rect 3997 1426 4074 1430
rect 3647 1421 3829 1424
rect 3447 1420 3829 1421
rect 3217 1418 3651 1420
rect 3011 1417 3651 1418
rect 3011 1416 3462 1417
rect 3011 1415 3228 1416
rect 4003 1414 4007 1426
rect 4051 1414 4055 1426
rect 3101 1399 3486 1401
rect 3101 1395 4004 1399
rect 4041 1394 4045 1408
rect 4059 1394 4063 1408
rect 4134 1394 4139 1606
rect 4271 1602 4275 1608
rect 4262 1598 4275 1602
rect 4262 1594 4266 1598
rect 4253 1583 4257 1590
rect 4271 1583 4275 1590
rect 4246 1579 4279 1583
rect 3350 1388 4014 1392
rect 4041 1390 4052 1394
rect 4059 1390 4139 1394
rect 4320 1505 4326 1644
rect 4390 1584 4396 1728
rect 4390 1552 4396 1579
rect 3583 1381 4024 1385
rect 2873 1286 2880 1380
rect 3881 1374 4033 1378
rect 4041 1370 4045 1390
rect 4012 1366 4045 1370
rect 4012 1362 4016 1366
rect 4031 1362 4035 1366
rect 4059 1362 4063 1390
rect 4003 1351 4007 1358
rect 4021 1351 4025 1358
rect 4041 1351 4045 1358
rect 4051 1351 4055 1358
rect 3836 1347 4074 1351
rect 4320 1307 4326 1499
rect 3068 1304 4327 1307
rect 3085 1298 3088 1304
rect 3141 1298 3144 1304
rect 3338 1298 3341 1304
rect 3601 1298 3604 1304
rect 2873 1283 3081 1286
rect 2875 1282 3081 1283
rect 3092 1285 3095 1294
rect 3092 1282 3099 1285
rect 3092 1278 3095 1282
rect 3128 1282 3137 1286
rect 3148 1285 3151 1294
rect 3148 1282 3165 1285
rect 3314 1282 3334 1286
rect 3345 1285 3348 1294
rect 3345 1282 3370 1285
rect 3148 1278 3151 1282
rect 3345 1278 3348 1282
rect 3572 1282 3597 1286
rect 3608 1285 3611 1294
rect 3608 1282 3707 1285
rect 3608 1278 3611 1282
rect 3085 1270 3088 1274
rect 3141 1270 3144 1274
rect 3338 1270 3341 1274
rect 3601 1270 3604 1274
rect 4390 1270 4396 1546
rect 3084 1267 3829 1270
rect 3099 1266 3103 1267
rect 3836 1267 4396 1270
rect 4442 1171 4448 1799
rect 2486 1170 4448 1171
rect 1760 1167 4448 1170
rect 1766 1152 1770 1167
rect 1785 1152 1789 1167
rect 1809 1152 1813 1167
rect 1852 1152 1856 1167
rect 1871 1152 1875 1167
rect 1895 1152 1899 1167
rect 1942 1152 1946 1167
rect 1961 1152 1965 1167
rect 1985 1152 1989 1167
rect 2037 1152 2041 1167
rect 2056 1152 2060 1167
rect 2080 1152 2084 1167
rect 2121 1152 2125 1167
rect 2140 1152 2144 1167
rect 2164 1152 2168 1167
rect 2207 1152 2211 1167
rect 2226 1152 2230 1167
rect 2250 1152 2254 1167
rect 2297 1152 2301 1167
rect 2316 1152 2320 1167
rect 2340 1152 2344 1167
rect 2392 1152 2396 1167
rect 2411 1152 2415 1167
rect 2435 1152 2439 1167
rect 2486 1166 4448 1167
rect 1775 1138 1779 1146
rect 1685 1134 1767 1138
rect 1775 1134 1810 1138
rect 1755 1125 1777 1129
rect 1785 1120 1789 1134
rect 1817 1120 1821 1146
rect 1861 1138 1865 1146
rect 1826 1134 1830 1138
rect 1841 1133 1845 1138
rect 1850 1134 1853 1138
rect 1861 1134 1896 1138
rect 1840 1125 1863 1129
rect 1871 1120 1875 1134
rect 1903 1120 1907 1146
rect 1951 1138 1955 1146
rect 1993 1138 1997 1146
rect 2046 1138 2050 1146
rect 2088 1138 2092 1146
rect 2130 1138 2134 1146
rect 2172 1138 2176 1146
rect 2216 1138 2220 1146
rect 2258 1138 2262 1146
rect 2306 1138 2310 1146
rect 2348 1138 2352 1146
rect 2401 1138 2405 1146
rect 2443 1138 2447 1146
rect 1912 1134 1916 1138
rect 1931 1134 1935 1138
rect 1940 1134 1943 1138
rect 1951 1134 1986 1138
rect 1993 1134 2001 1138
rect 1930 1125 1953 1129
rect 1961 1120 1965 1134
rect 1993 1120 1997 1134
rect 2026 1134 2030 1138
rect 2035 1134 2038 1138
rect 2046 1134 2081 1138
rect 2088 1134 2095 1138
rect 2024 1125 2048 1129
rect 2056 1120 2060 1134
rect 2088 1120 2092 1134
rect 2100 1134 2101 1138
rect 2110 1134 2114 1138
rect 2119 1134 2122 1138
rect 2130 1134 2165 1138
rect 2172 1134 2179 1138
rect 2110 1125 2132 1129
rect 2140 1120 2144 1134
rect 2172 1120 2176 1134
rect 2196 1134 2200 1138
rect 2205 1134 2208 1138
rect 2216 1134 2251 1138
rect 2258 1134 2267 1138
rect 2195 1125 2218 1129
rect 2226 1120 2230 1134
rect 2258 1120 2262 1134
rect 2286 1134 2290 1138
rect 2295 1134 2298 1138
rect 2306 1134 2341 1138
rect 2348 1134 2356 1138
rect 2285 1125 2308 1129
rect 2316 1120 2320 1134
rect 2348 1120 2352 1134
rect 2381 1134 2385 1138
rect 2390 1134 2393 1138
rect 2401 1134 2436 1138
rect 2443 1134 2452 1138
rect 2379 1125 2403 1129
rect 2411 1120 2415 1134
rect 2443 1120 2447 1134
rect 1766 1109 1770 1116
rect 1809 1109 1813 1116
rect 1852 1109 1856 1116
rect 1895 1109 1899 1116
rect 1942 1109 1946 1116
rect 1985 1109 1989 1116
rect 2037 1109 2041 1116
rect 2080 1109 2084 1116
rect 2121 1109 2125 1116
rect 2164 1109 2168 1116
rect 2207 1109 2211 1116
rect 2250 1109 2254 1116
rect 2297 1109 2301 1116
rect 2340 1109 2344 1116
rect 2392 1109 2396 1116
rect 2435 1109 2439 1116
rect 1759 1106 2450 1109
rect 1801 1094 1853 1099
rect 2019 1081 2024 1098
rect 2212 1087 2286 1092
rect 2212 1083 2217 1087
rect 1920 1078 2024 1081
rect 2091 1078 2217 1083
rect 1154 1069 1831 1070
rect 2486 1069 2490 1166
rect 2516 1165 4448 1166
rect 1154 1066 2492 1069
rect 1828 1051 1832 1066
rect 1847 1051 1851 1066
rect 1871 1051 1875 1066
rect 1914 1051 1918 1066
rect 1933 1051 1937 1066
rect 1957 1051 1961 1066
rect 2004 1051 2008 1066
rect 2023 1051 2027 1066
rect 2047 1051 2051 1066
rect 2099 1051 2103 1066
rect 2118 1051 2122 1066
rect 2142 1051 2146 1066
rect 1837 1037 1841 1045
rect 1879 1037 1883 1045
rect 1923 1037 1927 1045
rect 1965 1037 1969 1045
rect 1818 1033 1821 1037
rect 1826 1033 1829 1037
rect 1837 1033 1872 1037
rect 1879 1033 1892 1037
rect 1903 1033 1905 1037
rect 1801 1024 1839 1028
rect 1847 1019 1851 1033
rect 1879 1019 1883 1033
rect 1910 1033 1915 1037
rect 1923 1033 1958 1037
rect 1965 1033 1978 1037
rect 2013 1037 2017 1045
rect 2055 1037 2059 1045
rect 1996 1033 2005 1037
rect 2013 1033 2048 1037
rect 2055 1033 2068 1037
rect 2108 1037 2112 1045
rect 2150 1037 2154 1045
rect 2090 1033 2100 1037
rect 2108 1033 2143 1037
rect 2150 1033 2163 1037
rect 1903 1024 1910 1028
rect 1915 1024 1925 1028
rect 1933 1019 1937 1033
rect 1965 1019 1969 1033
rect 1997 1024 2015 1028
rect 2023 1019 2027 1033
rect 2055 1019 2059 1033
rect 2091 1024 2110 1028
rect 2118 1019 2122 1033
rect 2150 1019 2154 1033
rect 1828 1008 1832 1015
rect 1871 1008 1875 1015
rect 1914 1008 1918 1015
rect 1957 1008 1961 1015
rect 2004 1008 2008 1015
rect 2047 1008 2051 1015
rect 2099 1008 2103 1015
rect 2142 1008 2146 1015
rect 1127 1005 2156 1008
rect 1127 1004 1831 1005
rect 2267 995 2273 1020
rect 1997 990 2273 995
rect 2501 961 2507 1133
rect 2090 957 2507 961
rect 2090 956 2505 957
<< m2contact >>
rect 1646 3381 1651 3386
rect 1605 3365 1610 3370
rect 1808 3390 1813 3395
rect 1707 3381 1712 3386
rect 1725 3372 1732 3378
rect 1687 3365 1692 3370
rect 1754 3372 1760 3378
rect 1767 3374 1772 3379
rect 1869 3390 1874 3395
rect 1987 3392 1992 3397
rect 2045 3400 2050 3405
rect 1849 3374 1854 3379
rect 2004 3384 2009 3389
rect 2152 3400 2157 3405
rect 2086 3384 2091 3389
rect 1864 3266 1872 3273
rect 1987 3269 1992 3274
rect 1966 3196 1974 3202
rect 2058 3196 2065 3202
rect 2120 3200 2125 3205
rect 2113 3170 2120 3175
rect 2154 3200 2159 3205
rect 2129 3102 2134 3107
rect 1655 3049 1660 3054
rect 1614 3033 1619 3038
rect 1817 3058 1822 3063
rect 1716 3049 1721 3054
rect 1734 3040 1741 3046
rect 1696 3033 1701 3038
rect 1763 3040 1769 3046
rect 1776 3042 1781 3047
rect 1878 3058 1883 3063
rect 1996 3060 2001 3065
rect 2054 3068 2059 3073
rect 1858 3042 1863 3047
rect 2013 3052 2018 3057
rect 2161 3068 2166 3073
rect 2095 3052 2100 3057
rect 1873 2934 1881 2941
rect 1996 2937 2001 2942
rect 1975 2864 1983 2870
rect 2067 2864 2074 2870
rect 2129 2868 2134 2873
rect 2163 2868 2168 2873
rect 2293 3116 2301 3121
rect 2145 2745 2150 2750
rect 1676 2683 1681 2688
rect 1211 2525 1218 2532
rect 1635 2667 1640 2672
rect 1838 2692 1843 2697
rect 1737 2683 1742 2688
rect 1717 2667 1722 2672
rect 1755 2674 1762 2680
rect 1784 2674 1790 2680
rect 1797 2676 1802 2681
rect 1899 2692 1904 2697
rect 2017 2694 2022 2699
rect 2075 2702 2080 2707
rect 1879 2676 1884 2681
rect 2034 2686 2039 2691
rect 2182 2702 2187 2707
rect 2116 2686 2121 2691
rect 1894 2568 1902 2575
rect 1737 2525 1743 2530
rect 2017 2571 2022 2576
rect 1996 2498 2004 2504
rect 2088 2498 2095 2504
rect 2150 2502 2155 2507
rect 2184 2502 2189 2507
rect 2173 2362 2178 2368
rect 1704 2309 1709 2314
rect 1261 2292 1267 2297
rect 1663 2293 1668 2298
rect 1866 2318 1871 2323
rect 1765 2309 1770 2314
rect 1745 2293 1750 2298
rect 1783 2300 1790 2306
rect 1812 2300 1818 2306
rect 1825 2302 1830 2307
rect 1927 2318 1932 2323
rect 2045 2320 2050 2325
rect 2103 2328 2108 2333
rect 1907 2302 1912 2307
rect 2062 2312 2067 2317
rect 2210 2328 2215 2333
rect 2144 2312 2149 2317
rect 1922 2194 1930 2201
rect 2045 2197 2050 2202
rect 2024 2124 2032 2130
rect 2116 2124 2123 2130
rect 2178 2128 2183 2133
rect 2168 2098 2176 2103
rect 2212 2128 2217 2133
rect 2293 2745 2301 2750
rect 2293 2378 2301 2383
rect 2248 2098 2255 2103
rect 2525 2098 2533 2107
rect 2157 1908 2164 1913
rect 2471 1812 2478 1819
rect 2379 1789 2386 1797
rect 2736 1854 2744 1862
rect 1148 1733 1153 1738
rect 1063 1710 1068 1715
rect 1090 1710 1095 1716
rect 1119 1693 1124 1699
rect 1148 1667 1153 1672
rect 963 1634 968 1639
rect 1119 1605 1124 1610
rect 1148 1582 1153 1587
rect 1727 1739 1733 1744
rect 1704 1695 1710 1700
rect 1727 1685 1733 1690
rect 1812 1686 1818 1691
rect 1902 1686 1908 1691
rect 1997 1685 2002 1690
rect 2082 1685 2088 1690
rect 2167 1686 2173 1691
rect 2257 1686 2263 1691
rect 2352 1685 2357 1690
rect 2429 1665 2434 1670
rect 1261 1549 1266 1554
rect 1133 1527 1139 1533
rect 1119 1520 1124 1525
rect 1148 1493 1153 1498
rect 1705 1495 1711 1500
rect 963 1460 968 1465
rect 975 1451 980 1456
rect 1680 1451 1686 1456
rect 1705 1441 1711 1446
rect 1781 1450 1786 1455
rect 1790 1442 1796 1447
rect 1867 1450 1872 1455
rect 1880 1442 1886 1447
rect 1958 1450 1963 1455
rect 1975 1441 1980 1446
rect 2051 1450 2056 1455
rect 2060 1441 2066 1446
rect 2135 1450 2140 1455
rect 2145 1442 2151 1447
rect 2221 1450 2226 1455
rect 2235 1442 2241 1447
rect 2311 1450 2316 1455
rect 2330 1441 2335 1446
rect 1119 1431 1124 1436
rect 2405 1421 2412 1426
rect 1148 1410 1154 1415
rect 1781 1408 1786 1413
rect 1867 1380 1872 1385
rect 975 1368 980 1373
rect 1119 1349 1124 1354
rect 1958 1356 1963 1361
rect 2051 1343 2056 1348
rect 2135 1320 2140 1325
rect 2221 1301 2226 1306
rect 2311 1291 2316 1296
rect 1749 1178 1755 1183
rect 2795 1788 2803 1797
rect 3144 1768 3151 1773
rect 3393 1761 3399 1766
rect 3637 1753 3644 1759
rect 3820 1674 3825 1679
rect 2994 1640 2999 1645
rect 2953 1624 2958 1629
rect 3055 1640 3060 1645
rect 3144 1639 3149 1644
rect 3243 1640 3248 1645
rect 3035 1624 3040 1629
rect 3202 1624 3207 1629
rect 3304 1640 3309 1645
rect 3393 1639 3398 1644
rect 3500 1640 3505 1645
rect 3284 1624 3289 1629
rect 3459 1624 3464 1629
rect 3561 1640 3566 1645
rect 3637 1639 3642 1644
rect 3722 1640 3727 1645
rect 3541 1624 3546 1629
rect 3657 1631 3663 1636
rect 3671 1623 3677 1628
rect 3681 1624 3686 1629
rect 3783 1640 3788 1645
rect 4028 1729 4034 1734
rect 3763 1624 3768 1629
rect 4319 1674 4326 1681
rect 3841 1547 3847 1552
rect 3307 1521 3316 1532
rect 3598 1522 3606 1529
rect 3826 1500 3833 1506
rect 4068 1500 4075 1505
rect 3143 1461 3150 1467
rect 3417 1456 3423 1462
rect 3598 1466 3604 1472
rect 2986 1433 2992 1439
rect 3095 1442 3100 1447
rect 3165 1439 3172 1447
rect 3344 1447 3350 1452
rect 3432 1447 3440 1454
rect 3370 1434 3375 1439
rect 3576 1456 3583 1461
rect 3626 1458 3633 1464
rect 3644 1452 3650 1457
rect 3657 1444 3665 1450
rect 3730 1431 3736 1436
rect 3874 1466 3881 1471
rect 3095 1395 3101 1401
rect 4279 1579 4284 1584
rect 3344 1387 3350 1392
rect 4390 1728 4397 1734
rect 4390 1579 4399 1584
rect 4390 1546 4397 1552
rect 4320 1499 4327 1505
rect 3576 1380 3583 1385
rect 3874 1373 3881 1378
rect 3099 1281 3104 1286
rect 3165 1282 3170 1287
rect 3370 1281 3375 1286
rect 3566 1282 3572 1287
rect 3707 1282 3712 1287
rect 3077 1265 3084 1270
rect 1680 1134 1685 1139
rect 1749 1124 1755 1129
rect 1821 1133 1826 1138
rect 1834 1125 1840 1130
rect 1907 1133 1912 1138
rect 1924 1125 1930 1130
rect 2001 1133 2006 1138
rect 2019 1124 2024 1129
rect 2095 1133 2100 1138
rect 2104 1124 2110 1129
rect 2179 1133 2185 1138
rect 2189 1125 2195 1130
rect 2267 1133 2272 1138
rect 2279 1125 2285 1130
rect 2356 1133 2362 1138
rect 2374 1124 2379 1129
rect 2452 1133 2458 1138
rect 2450 1105 2455 1110
rect 1796 1094 1801 1099
rect 1853 1094 1858 1099
rect 2019 1098 2024 1103
rect 1915 1077 1920 1082
rect 2286 1087 2291 1092
rect 2084 1077 2091 1083
rect 1146 1065 1154 1070
rect 2501 1133 2507 1138
rect 1821 1032 1826 1037
rect 1796 1023 1801 1028
rect 1905 1032 1910 1037
rect 1991 1033 1996 1038
rect 2084 1033 2090 1038
rect 1910 1023 1915 1028
rect 1991 1023 1997 1028
rect 2085 1023 2091 1028
rect 2267 1020 2273 1025
rect 1119 1004 1127 1009
rect 2156 1005 2163 1010
rect 1991 990 1997 995
rect 2083 956 2090 961
<< metal2 >>
rect 1367 3663 2476 3667
rect 1367 3029 1371 3663
rect 1725 3547 1732 3548
rect 1725 3540 2405 3547
rect 1651 3381 1707 3385
rect 1725 3378 1732 3540
rect 2050 3400 2152 3404
rect 1813 3390 1869 3394
rect 1732 3372 1754 3378
rect 1772 3374 1849 3379
rect 1610 3365 1687 3370
rect 1754 3273 1760 3372
rect 1987 3274 1992 3392
rect 2009 3384 2086 3389
rect 1754 3266 1864 3273
rect 1987 3268 1992 3269
rect 1974 3196 2058 3202
rect 2125 3200 2154 3204
rect 2120 3170 2248 3175
rect 2263 3138 2333 3144
rect 1734 3129 1741 3132
rect 2263 3129 2269 3138
rect 1734 3123 2269 3129
rect 1660 3049 1716 3053
rect 1734 3046 1741 3123
rect 2129 3116 2293 3119
rect 2129 3107 2134 3116
rect 2059 3068 2161 3072
rect 1822 3058 1878 3062
rect 1741 3040 1763 3046
rect 1781 3042 1858 3047
rect 1619 3033 1696 3038
rect 1614 3029 1619 3033
rect 1367 3025 1619 3029
rect 1763 2941 1769 3040
rect 1996 2942 2001 3060
rect 2018 3052 2095 3057
rect 1763 2934 1873 2941
rect 1996 2936 2001 2937
rect 1983 2864 2067 2870
rect 2134 2868 2163 2872
rect 2121 2838 2248 2843
rect 2150 2745 2293 2750
rect 2080 2702 2182 2706
rect 1843 2692 1899 2696
rect 1681 2683 1737 2687
rect 1762 2674 1784 2680
rect 1802 2676 1879 2681
rect 1640 2667 1717 2672
rect 1784 2575 1790 2674
rect 2017 2576 2022 2694
rect 2039 2686 2116 2691
rect 1784 2568 1894 2575
rect 2017 2570 2022 2571
rect 1218 2525 1737 2530
rect 2004 2498 2088 2504
rect 2155 2502 2184 2506
rect 2141 2472 2248 2477
rect 2173 2378 2293 2382
rect 2173 2368 2178 2378
rect 2108 2328 2210 2332
rect 1871 2318 1927 2322
rect 1709 2309 1765 2313
rect 1790 2300 1812 2306
rect 1830 2302 1907 2307
rect 1668 2293 1745 2298
rect 1065 1691 1068 1710
rect 961 1688 1068 1691
rect 963 1639 967 1688
rect 1091 1683 1094 1710
rect 975 1680 1094 1683
rect 963 1465 967 1634
rect 975 1456 979 1680
rect 1119 1610 1124 1693
rect 1119 1533 1124 1605
rect 1148 1672 1153 1733
rect 1148 1587 1153 1667
rect 1119 1527 1133 1533
rect 1119 1525 1124 1527
rect 975 1373 979 1451
rect 1119 1436 1124 1520
rect 1119 1357 1124 1431
rect 1148 1498 1153 1582
rect 1261 1554 1266 2292
rect 1812 2201 1818 2300
rect 2045 2202 2050 2320
rect 2067 2312 2144 2317
rect 1812 2194 1922 2201
rect 2045 2196 2050 2197
rect 2032 2124 2116 2130
rect 2183 2128 2212 2132
rect 2176 2098 2248 2103
rect 2328 1912 2332 3138
rect 2164 1908 2332 1912
rect 2398 1798 2405 3540
rect 2472 1862 2476 3663
rect 2526 2107 2532 2109
rect 2471 1819 2477 1862
rect 2379 1797 2405 1798
rect 2386 1791 2405 1797
rect 2526 1764 2532 2098
rect 2744 1854 3677 1861
rect 2803 1791 3663 1797
rect 1733 1739 2357 1744
rect 1704 1525 1710 1695
rect 1727 1690 1733 1739
rect 1812 1691 1818 1739
rect 1902 1691 1908 1739
rect 1997 1690 2002 1739
rect 2082 1690 2088 1739
rect 2167 1691 2173 1739
rect 2257 1691 2263 1739
rect 2352 1690 2357 1739
rect 2525 1670 2533 1764
rect 2434 1665 2533 1670
rect 1148 1421 1153 1493
rect 1147 1415 1153 1421
rect 1680 1521 1710 1525
rect 1680 1461 1684 1521
rect 1711 1495 2335 1500
rect 1680 1456 1685 1461
rect 1147 1410 1148 1415
rect 1119 1354 1125 1357
rect 1124 1349 1125 1354
rect 1119 1050 1125 1349
rect 1147 1112 1153 1410
rect 1680 1139 1685 1451
rect 1705 1446 1711 1495
rect 1781 1413 1786 1450
rect 1790 1447 1796 1495
rect 1867 1385 1872 1450
rect 1880 1447 1886 1495
rect 1958 1361 1963 1450
rect 1975 1446 1980 1495
rect 2051 1348 2056 1450
rect 2060 1446 2066 1495
rect 2135 1325 2140 1450
rect 2145 1447 2151 1495
rect 2221 1306 2226 1450
rect 2235 1447 2241 1495
rect 2311 1296 2316 1450
rect 2330 1446 2335 1495
rect 2525 1426 2533 1665
rect 2999 1640 3055 1644
rect 3144 1644 3149 1768
rect 3248 1640 3304 1644
rect 3393 1644 3398 1761
rect 2958 1624 3035 1629
rect 3144 1532 3149 1639
rect 3505 1640 3561 1644
rect 3637 1644 3642 1753
rect 3642 1639 3650 1643
rect 3207 1624 3284 1629
rect 3393 1553 3398 1639
rect 3464 1624 3541 1629
rect 3393 1547 3633 1553
rect 3144 1528 3307 1532
rect 3144 1467 3149 1528
rect 3393 1523 3398 1547
rect 3308 1471 3314 1521
rect 3393 1518 3439 1523
rect 3308 1467 3423 1471
rect 3418 1462 3423 1467
rect 3432 1454 3440 1518
rect 3598 1472 3604 1522
rect 3626 1464 3633 1547
rect 2412 1421 2533 1426
rect 2525 1270 2533 1421
rect 2986 1365 2992 1433
rect 3095 1401 3100 1442
rect 2986 1362 3115 1365
rect 3112 1285 3115 1362
rect 3166 1287 3170 1439
rect 3344 1392 3350 1447
rect 3104 1282 3115 1285
rect 3370 1286 3375 1434
rect 3576 1385 3583 1456
rect 3644 1457 3650 1639
rect 3657 1636 3663 1791
rect 3657 1450 3663 1631
rect 3671 1628 3677 1854
rect 4034 1729 4390 1734
rect 3825 1674 4319 1679
rect 3727 1640 3783 1644
rect 3686 1624 3763 1629
rect 3671 1356 3677 1623
rect 4284 1579 4390 1584
rect 3847 1547 4390 1552
rect 3833 1500 4068 1504
rect 4075 1500 4320 1504
rect 3707 1431 3730 1436
rect 3671 1351 3678 1356
rect 3566 1345 3678 1351
rect 3566 1287 3572 1345
rect 3707 1287 3712 1431
rect 3874 1378 3881 1466
rect 2524 1265 3077 1270
rect 1755 1178 2379 1183
rect 1749 1129 1755 1178
rect 1147 1070 1154 1112
rect 1119 1009 1126 1050
rect 1796 1028 1801 1094
rect 1821 1037 1826 1133
rect 1834 1130 1840 1178
rect 1907 1098 1912 1133
rect 1924 1130 1930 1178
rect 1858 1094 1912 1098
rect 2001 1090 2006 1133
rect 2019 1129 2024 1178
rect 2095 1102 2100 1133
rect 2104 1129 2110 1178
rect 2024 1098 2100 1102
rect 2179 1093 2185 1133
rect 2189 1130 2195 1178
rect 1905 1087 2006 1090
rect 2013 1089 2185 1093
rect 1905 1037 1910 1087
rect 1915 1024 1920 1077
rect 2013 1075 2017 1089
rect 1991 1072 2017 1075
rect 1991 1038 1996 1072
rect 2085 1038 2089 1077
rect 1991 995 1997 1023
rect 2085 961 2091 1023
rect 2267 1025 2272 1133
rect 2279 1130 2285 1178
rect 2356 1092 2362 1133
rect 2374 1129 2379 1178
rect 2458 1133 2501 1138
rect 2525 1114 2533 1265
rect 2524 1110 2533 1114
rect 2455 1105 2533 1110
rect 2291 1087 2362 1092
rect 2267 1019 2272 1020
rect 2524 1010 2533 1105
rect 2163 1005 2534 1010
rect 2090 956 2091 961
<< m123contact >>
rect 2135 3433 2141 3438
rect 1581 3364 1586 3369
rect 1691 3331 1697 3336
rect 1724 3330 1732 3336
rect 1864 3341 1869 3347
rect 1768 3330 1773 3336
rect 1957 3310 1962 3315
rect 2005 3350 2010 3356
rect 2016 3310 2024 3315
rect 2112 3310 2120 3315
rect 2135 3311 2143 3316
rect 1864 3249 1869 3254
rect 1956 3249 1961 3254
rect 2019 3249 2024 3254
rect 2112 3235 2120 3241
rect 2054 3170 2064 3175
rect 2248 3170 2255 3175
rect 2159 3142 2164 3147
rect 2144 3101 2150 3106
rect 1703 3000 1708 3005
rect 1733 2998 1741 3004
rect 1873 3009 1878 3015
rect 1777 2998 1782 3004
rect 1966 2978 1971 2983
rect 2014 3019 2019 3024
rect 2025 2978 2033 2983
rect 2121 2978 2129 2983
rect 2144 2979 2151 2984
rect 1873 2917 1878 2922
rect 1965 2917 1970 2922
rect 2028 2917 2033 2922
rect 2121 2903 2129 2909
rect 2063 2838 2073 2843
rect 2248 2838 2256 2843
rect 2166 2773 2173 2781
rect 2165 2735 2171 2740
rect 1626 2666 1631 2671
rect 1722 2633 1728 2639
rect 1754 2632 1762 2638
rect 1894 2643 1899 2649
rect 1798 2632 1803 2638
rect 1987 2612 1992 2617
rect 2035 2653 2040 2658
rect 2046 2612 2054 2617
rect 2142 2612 2150 2617
rect 2165 2613 2172 2618
rect 1894 2551 1899 2557
rect 1986 2551 1991 2556
rect 2049 2551 2054 2556
rect 2142 2537 2150 2543
rect 2084 2472 2094 2477
rect 2248 2472 2254 2478
rect 2188 2405 2194 2411
rect 2193 2360 2199 2366
rect 1602 2306 1607 2311
rect 1127 1710 1132 1715
rect 988 1625 993 1630
rect 988 1540 993 1545
rect 1750 2259 1755 2264
rect 1782 2258 1790 2264
rect 1922 2269 1927 2275
rect 1826 2258 1831 2264
rect 2015 2238 2020 2243
rect 2063 2279 2068 2284
rect 2074 2238 2082 2243
rect 2170 2238 2178 2243
rect 2193 2239 2200 2245
rect 1922 2177 1928 2182
rect 2014 2177 2020 2182
rect 2077 2177 2082 2182
rect 2170 2163 2178 2169
rect 1799 2093 1804 2099
rect 2112 2098 2122 2103
rect 2243 1812 2250 1819
rect 1563 1799 1569 1804
rect 2073 1799 2078 1804
rect 1983 1785 1988 1790
rect 2157 1786 2163 1792
rect 2333 1789 2340 1797
rect 2666 1811 2675 1824
rect 1799 1694 1804 1699
rect 1823 1694 1828 1699
rect 1890 1694 1895 1699
rect 1913 1694 1918 1699
rect 1983 1694 1988 1699
rect 2008 1694 2013 1699
rect 2073 1694 2078 1699
rect 2092 1694 2097 1699
rect 2157 1694 2162 1699
rect 2178 1694 2183 1699
rect 2243 1694 2248 1699
rect 2268 1694 2273 1699
rect 2334 1694 2339 1699
rect 2363 1694 2368 1699
rect 2429 1694 2434 1699
rect 2709 1742 2720 1754
rect 2641 1715 2651 1725
rect 2940 1687 2950 1696
rect 1801 1450 1806 1455
rect 1891 1450 1896 1455
rect 1986 1450 1991 1455
rect 2070 1450 2075 1455
rect 2156 1450 2161 1455
rect 2246 1450 2251 1455
rect 2341 1450 2346 1455
rect 2407 1450 2412 1455
rect 2940 1622 2946 1628
rect 3162 1631 3167 1636
rect 3171 1622 3177 1628
rect 3437 1631 3443 1636
rect 3412 1624 3419 1629
rect 2795 1450 2803 1456
rect 2434 1408 2441 1413
rect 2434 1380 2440 1385
rect 2436 1356 2444 1361
rect 2436 1343 2446 1348
rect 2436 1320 2445 1325
rect 2438 1300 2445 1306
rect 2454 1291 2460 1296
rect 2917 1408 2925 1414
rect 2873 1380 2880 1385
rect 2641 1343 2650 1349
rect 2667 1319 2675 1326
rect 2710 1300 2720 1307
rect 2737 1291 2744 1296
rect 3185 1431 3190 1436
rect 3123 1281 3128 1286
rect 3309 1282 3314 1287
rect 3437 1426 3444 1431
rect 3829 1419 3836 1424
rect 3829 1345 3836 1351
rect 3829 1265 3836 1270
rect 1845 1133 1850 1138
rect 1935 1133 1940 1138
rect 2030 1133 2035 1138
rect 2114 1133 2119 1138
rect 2200 1133 2205 1138
rect 2290 1133 2295 1138
rect 2385 1133 2390 1138
<< metal3 >>
rect 1439 3578 2434 3583
rect 1439 3369 1444 3578
rect 1438 3364 1581 3369
rect 2005 3346 2010 3350
rect 1869 3342 2010 3346
rect 1691 3254 1697 3331
rect 1732 3330 1768 3336
rect 1864 3254 1869 3341
rect 2135 3316 2141 3433
rect 1962 3310 2016 3314
rect 1691 3249 1864 3254
rect 1961 3249 2019 3252
rect 1992 3175 1996 3249
rect 2112 3241 2119 3310
rect 1992 3170 2054 3175
rect 1740 3142 2159 3147
rect 1741 3004 1747 3142
rect 2014 3014 2019 3019
rect 1878 3010 2019 3014
rect 1703 2922 1708 3000
rect 1741 2998 1777 3004
rect 1873 2922 1878 3009
rect 2144 2984 2150 3101
rect 1971 2978 2025 2982
rect 1703 2917 1873 2922
rect 1970 2917 2028 2920
rect 1703 2915 1708 2917
rect 2001 2843 2005 2917
rect 2121 2909 2128 2978
rect 2001 2838 2063 2843
rect 1762 2773 2166 2781
rect 1563 2666 1626 2671
rect 1563 1804 1568 2666
rect 1763 2638 1769 2773
rect 2035 2648 2040 2653
rect 1899 2644 2040 2648
rect 1722 2556 1728 2633
rect 1762 2632 1798 2638
rect 1894 2557 1899 2643
rect 2165 2618 2171 2735
rect 1992 2612 2046 2616
rect 1722 2551 1894 2556
rect 1991 2551 2049 2554
rect 2022 2477 2026 2551
rect 2142 2543 2149 2612
rect 2022 2472 2084 2477
rect 1800 2405 2188 2411
rect 1602 2131 1607 2306
rect 1800 2264 1807 2405
rect 2063 2274 2068 2279
rect 1927 2270 2068 2274
rect 1750 2182 1755 2259
rect 1790 2258 1826 2264
rect 1922 2182 1927 2269
rect 2193 2245 2199 2360
rect 2020 2238 2074 2242
rect 1750 2177 1922 2182
rect 2020 2177 2077 2180
rect 1602 2127 1895 2131
rect 1128 1678 1132 1710
rect 1799 1699 1804 2093
rect 1890 1699 1895 2127
rect 2050 2103 2054 2177
rect 2170 2169 2177 2238
rect 2050 2098 2112 2103
rect 1983 1699 1988 1785
rect 2073 1699 2078 1799
rect 2157 1699 2162 1786
rect 2243 1699 2248 1812
rect 2334 1699 2339 1789
rect 2429 1699 2434 3578
rect 2675 1819 3443 1824
rect 2675 1818 2862 1819
rect 2720 1753 2812 1754
rect 2720 1748 3418 1753
rect 2720 1747 2812 1748
rect 2769 1725 3131 1726
rect 2651 1718 3131 1725
rect 2651 1717 2796 1718
rect 3123 1697 3130 1718
rect 988 1675 1132 1678
rect 988 1630 993 1675
rect 1823 1637 1828 1694
rect 988 1545 993 1625
rect 1801 1633 1828 1637
rect 1801 1455 1806 1633
rect 1913 1588 1918 1694
rect 2008 1624 2013 1694
rect 2092 1624 2097 1694
rect 2178 1624 2183 1694
rect 2268 1626 2273 1694
rect 1986 1621 2013 1624
rect 2070 1621 2097 1624
rect 2156 1621 2183 1624
rect 2246 1623 2273 1626
rect 2363 1625 2368 1694
rect 1801 1396 1806 1450
rect 1891 1585 1919 1588
rect 1891 1455 1896 1585
rect 1801 1393 1849 1396
rect 1801 1392 1806 1393
rect 1845 1138 1849 1393
rect 1891 1381 1896 1450
rect 1986 1455 1991 1621
rect 1986 1382 1991 1450
rect 2070 1455 2075 1621
rect 2070 1382 2075 1450
rect 2156 1455 2161 1621
rect 1891 1378 1940 1381
rect 1986 1379 2036 1382
rect 2070 1379 2119 1382
rect 1935 1138 1940 1378
rect 2031 1208 2036 1379
rect 2030 1169 2036 1208
rect 2030 1138 2035 1169
rect 2114 1138 2119 1379
rect 2156 1380 2161 1450
rect 2246 1455 2251 1623
rect 2200 1380 2205 1381
rect 2156 1377 2205 1380
rect 2200 1138 2205 1377
rect 2246 1379 2251 1450
rect 2341 1622 2368 1625
rect 3123 1692 3177 1697
rect 2940 1628 2946 1687
rect 2341 1455 2346 1622
rect 2412 1450 2795 1455
rect 2341 1380 2346 1450
rect 2441 1408 2917 1413
rect 2385 1380 2390 1381
rect 2440 1380 2873 1385
rect 2246 1376 2295 1379
rect 2341 1377 2390 1380
rect 2290 1138 2295 1376
rect 2385 1138 2390 1377
rect 2444 1356 2763 1361
rect 2446 1343 2641 1348
rect 2445 1320 2667 1325
rect 2675 1320 2676 1325
rect 2445 1300 2710 1306
rect 2720 1300 2721 1306
rect 2460 1291 2737 1296
rect 2756 1220 2763 1356
rect 3123 1286 3128 1692
rect 3162 1509 3166 1631
rect 3171 1628 3177 1692
rect 3413 1629 3418 1748
rect 3437 1636 3443 1819
rect 3162 1505 3190 1509
rect 3185 1436 3190 1505
rect 3185 1220 3190 1431
rect 3413 1428 3418 1624
rect 3309 1424 3418 1428
rect 3437 1431 3443 1631
rect 3309 1287 3314 1424
rect 3829 1351 3836 1419
rect 3829 1270 3836 1345
rect 2753 1212 3190 1220
<< labels >>
rlabel metal1 1097 1711 1101 1715 1 S1
rlabel metal1 1041 1711 1045 1715 3 S0
rlabel metal1 1042 1733 1123 1736 5 VDD
rlabel metal1 1042 1696 1123 1699 1 GND
rlabel metal1 1119 1711 1123 1714 7 S1not
rlabel metal1 1005 1667 1072 1670 1 VDD
rlabel metal1 1006 1582 1073 1585 1 VDD
rlabel metal1 1006 1493 1073 1496 1 VDD
rlabel metal1 1005 1521 1074 1524 1 GND
rlabel metal1 1005 1432 1074 1435 1 GND
rlabel metal1 1000 1625 1005 1629 3 S1not
rlabel metal1 1001 1549 1006 1553 3 S0
rlabel metal1 1001 1540 1006 1544 3 S1not
rlabel metal1 1001 1460 1006 1464 3 S0not
rlabel metal1 1001 1451 1006 1455 3 S1
rlabel metal1 1071 1634 1076 1638 1 D0
rlabel metal1 1072 1549 1077 1553 1 D1
rlabel metal1 1001 1368 1006 1372 3 S1
rlabel metal1 1001 1377 1006 1381 3 S0
rlabel metal1 1005 1349 1074 1352 1 GND
rlabel metal1 1006 1410 1073 1413 1 VDD
rlabel metal1 1072 1460 1077 1464 1 D2
rlabel metal1 1072 1377 1077 1381 1 D3
rlabel metal1 1004 1606 1073 1609 1 GND
rlabel m2contact 1063 1711 1067 1714 1 S0not
rlabel metal3 988 1675 993 1678 1 S1not
rlabel metal2 975 1680 979 1683 1 S1
rlabel metal2 961 1688 965 1691 1 S0not
rlabel metal1 955 1711 959 1715 3 S0
rlabel metal1 1000 1634 1005 1638 3 S0not
rlabel metal1 1734 1423 1744 1426 1 GND
rlabel metal1 1808 1423 1818 1426 1 GND
rlabel metal1 1891 1423 1901 1426 1 GND
rlabel metal1 1989 1423 1999 1426 1 GND
rlabel metal1 1738 1484 1748 1487 5 VDD
rlabel metal1 1806 1484 1816 1487 5 VDD
rlabel metal1 1903 1484 1913 1487 5 VDD
rlabel metal1 2001 1484 2011 1487 5 VDD
rlabel metal1 2089 1423 2099 1426 1 GND
rlabel metal1 2163 1423 2173 1426 1 GND
rlabel metal1 2246 1423 2256 1426 1 GND
rlabel metal1 2344 1423 2354 1426 1 GND
rlabel metal1 2093 1484 2103 1487 5 VDD
rlabel metal1 2161 1484 2171 1487 5 VDD
rlabel metal1 2258 1484 2268 1487 5 VDD
rlabel metal1 2356 1484 2366 1487 5 VDD
rlabel m2contact 1782 1451 1786 1455 1 compA3
rlabel metal1 2337 1451 2341 1455 1 B0
rlabel metal1 2400 1167 2410 1170 5 VDD
rlabel metal1 2302 1167 2312 1170 5 VDD
rlabel metal1 2205 1167 2215 1170 5 VDD
rlabel metal1 2137 1167 2147 1170 5 VDD
rlabel metal1 2388 1106 2398 1109 1 GND
rlabel metal1 2290 1106 2300 1109 1 GND
rlabel metal1 2207 1106 2217 1109 1 GND
rlabel metal1 2133 1106 2143 1109 1 GND
rlabel metal1 2045 1167 2055 1170 5 VDD
rlabel metal1 1947 1167 1957 1170 5 VDD
rlabel metal1 1850 1167 1860 1170 5 VDD
rlabel metal1 1782 1167 1792 1170 5 VDD
rlabel metal1 2033 1106 2043 1109 1 GND
rlabel metal1 1935 1106 1945 1109 1 GND
rlabel metal1 1852 1106 1862 1109 1 GND
rlabel metal1 1778 1106 1788 1109 1 GND
rlabel m2contact 2267 1134 2271 1138 1 AndB1
rlabel m2contact 2002 1134 2006 1138 1 AndA2
rlabel metal1 1840 1005 1850 1008 1 GND
rlabel metal1 1914 1005 1924 1008 1 GND
rlabel metal1 1997 1005 2007 1008 1 GND
rlabel metal1 2095 1005 2105 1008 1 GND
rlabel metal1 1844 1066 1854 1069 5 VDD
rlabel metal1 1912 1066 1922 1069 5 VDD
rlabel metal1 2009 1066 2019 1069 5 VDD
rlabel metal1 2107 1066 2117 1069 5 VDD
rlabel metal1 1743 1178 1749 1183 1 D3
rlabel metal1 1756 1667 1766 1670 1 GND
rlabel metal1 1830 1667 1840 1670 1 GND
rlabel metal1 1913 1667 1923 1670 1 GND
rlabel metal1 2011 1667 2021 1670 1 GND
rlabel metal1 1760 1728 1770 1731 5 VDD
rlabel metal1 1828 1728 1838 1731 5 VDD
rlabel metal1 1925 1728 1935 1731 5 VDD
rlabel metal1 2023 1728 2033 1731 5 VDD
rlabel metal1 2111 1667 2121 1670 1 GND
rlabel metal1 2185 1667 2195 1670 1 GND
rlabel metal1 2268 1667 2278 1670 1 GND
rlabel metal1 2366 1667 2376 1670 1 GND
rlabel metal1 2115 1728 2125 1731 5 VDD
rlabel metal1 2183 1728 2193 1731 5 VDD
rlabel metal1 2280 1728 2290 1731 5 VDD
rlabel metal1 2378 1728 2388 1731 5 VDD
rlabel metal1 1699 1495 1705 1500 1 D2
rlabel metal1 1888 1033 1892 1037 1 AndY3
rlabel metal1 1974 1033 1978 1037 1 AndY2
rlabel metal1 2064 1033 2068 1037 1 AndY1
rlabel metal1 2159 1033 2163 1037 1 AndY0
rlabel metal1 1551 1066 1559 1070 1 VDD
rlabel metal1 1556 1004 1564 1008 1 GND
rlabel metal1 1826 1134 1830 1138 1 AndA3
rlabel metal1 1912 1134 1916 1138 1 AndB3
rlabel metal1 1797 1451 1801 1455 1 B3
rlabel m2contact 1868 1451 1872 1455 1 CompB3
rlabel metal1 1841 1134 1845 1138 1 B3
rlabel metal1 1311 1593 1368 1598 5 VDD
rlabel metal1 1310 1527 1367 1532 1 GND
rlabel metal1 1225 1562 1229 1575 1 D0
rlabel metal1 1220 1549 1226 1553 1 D1
rlabel metal1 1721 1739 1727 1744 1 Eadd_sub
rlabel metal1 1804 1695 1808 1699 1 Add_subA3
rlabel metal1 1819 1695 1823 1699 1 B3
rlabel metal1 1909 1695 1913 1699 1 A2
rlabel metal1 1980 1695 1984 1699 1 Add_SubA2
rlabel metal1 2004 1695 2008 1699 1 B2
rlabel metal1 2075 1695 2079 1699 1 Add_SubB2
rlabel metal1 2088 1695 2092 1699 1 A1
rlabel metal1 2159 1695 2163 1699 1 Add_SubA1
rlabel metal1 2174 1695 2178 1699 1 B1
rlabel metal1 2245 1695 2249 1699 1 Add_SubB1
rlabel metal1 2264 1695 2268 1699 1 A0
rlabel metal1 2335 1695 2339 1699 1 Add_SubA0
rlabel metal1 2359 1695 2363 1699 1 B0
rlabel metal1 2429 1695 2433 1699 1 Add_SubB0
rlabel metal1 1714 1695 1718 1699 1 A3
rlabel metal1 1691 1451 1695 1455 1 A3
rlabel metal1 1690 1134 1694 1138 1 A3
rlabel metal1 1931 1134 1935 1138 1 A2
rlabel metal1 2026 1134 2030 1138 1 B2
rlabel metal1 2097 1134 2101 1138 1 AndB2
rlabel metal1 2110 1134 2114 1138 1 A1
rlabel m2contact 2181 1134 2185 1138 1 AndA1
rlabel metal1 2196 1134 2200 1138 1 B1
rlabel metal1 2286 1134 2290 1138 1 A0
rlabel m2contact 2357 1134 2361 1138 1 AndA0
rlabel metal1 2381 1134 2385 1138 1 B0
rlabel m2contact 2452 1134 2456 1138 1 AndB0
rlabel metal1 1887 1451 1891 1455 1 A2
rlabel m2contact 1958 1451 1962 1455 1 CompA2
rlabel metal1 1982 1451 1986 1455 1 B2
rlabel metal1 2053 1451 2057 1455 1 CompB2
rlabel metal1 2066 1451 2070 1455 1 A1
rlabel metal1 2137 1451 2141 1455 1 CompA1
rlabel metal1 2152 1451 2156 1455 1 B1
rlabel metal1 2223 1451 2227 1455 1 CompB1
rlabel metal1 2242 1451 2246 1455 1 A0
rlabel metal1 2313 1451 2317 1455 1 CompA0
rlabel metal1 2407 1451 2411 1455 1 CompB0
rlabel metal1 1818 1035 1820 1037 1 AndA3
rlabel metal1 1818 1026 1820 1028 1 AndB3
rlabel m2contact 2088 1035 2089 1037 1 AndA0
rlabel m2contact 2088 1026 2089 1028 1 AndB0
rlabel m2contact 1993 1026 1994 1028 1 AndB1
rlabel metal1 1903 1035 1904 1037 1 AndA2
rlabel metal1 1903 1026 1904 1028 1 AndB2
rlabel m2contact 1993 1035 1994 1037 1 AndA1
rlabel metal1 2217 2128 2222 2133 7 Carryout
rlabel metal1 2168 2868 2173 2873 1 Carry1
rlabel metal1 2189 2502 2194 2507 1 Carry2
rlabel metal1 1728 2998 1733 3004 1 Carry0
rlabel metal1 1777 2258 1782 2264 1 Carry2
rlabel metal1 1605 3415 1695 3419 1 VDD
rlabel metal1 1767 3424 1797 3428 1 VDD
rlabel metal1 2004 3434 2094 3438 5 VDD
rlabel metal1 1794 3092 1808 3096 1 VDD
rlabel metal1 2038 3102 2052 3106 1 VDD
rlabel metal1 2065 2979 2072 2982 1 VDD
rlabel metal1 1635 2717 1725 2721 1 VDD
rlabel metal1 2034 2736 2124 2740 5 VDD
rlabel metal1 1797 2726 1827 2730 1 VDD
rlabel metal1 1663 2343 1753 2347 1 VDD
rlabel metal1 1825 2352 1855 2356 1 VDD
rlabel metal1 2062 2362 2152 2366 5 VDD
rlabel metal1 1768 3341 1858 3345 1 GND
rlabel metal1 1783 3009 1797 3013 1 GND
rlabel metal1 2044 3019 2058 3023 1 GND
rlabel metal1 2060 2918 2067 2921 1 GND
rlabel metal1 1798 2643 1888 2647 1 GND
rlabel metal1 1640 3333 1642 3336 1 GND
rlabel metal1 1637 3084 1643 3087 1 VDD
rlabel metal1 1644 3000 1650 3003 1 GND
rlabel metal1 1875 2270 1882 2273 1 GND
rlabel metal1 2099 2279 2106 2282 1 GND
rlabel metal1 2293 3311 2301 3325 7 VDD
rlabel metal1 2248 2904 2254 2912 1 GND
rlabel metal1 1777 2300 1783 2306 1 Add_SubA3
rlabel metal1 1655 2301 1659 2305 1 Add_SubB3
rlabel metal1 1599 3374 1601 3376 1 D1
rlabel metal1 1588 3042 1590 3044 1 D1
rlabel metal1 1585 2676 1587 2678 1 D1
rlabel metal1 1570 2294 1572 2296 1 D1
rlabel metal1 1719 3330 1724 3336 1 D1
rlabel metal1 1597 3365 1603 3369 1 Add_SubB0
rlabel metal1 1719 3372 1725 3378 1 Add_SubA0
rlabel metal1 2215 2328 2221 2333 1 Add_SubS3
rlabel metal1 2187 2702 2193 2707 1 Add_SubS2
rlabel metal1 2166 3068 2172 3073 1 Add_SubS1
rlabel metal1 2157 3400 2163 3405 1 Add_SubS0
rlabel metal1 1606 3033 1611 3037 1 Add_SubB1
rlabel metal1 1728 3040 1734 3046 1 Add_SubA1
rlabel metal1 1627 2667 1631 2671 1 Add_SubB2
rlabel metal1 1749 2674 1755 2680 1 Add_SubA2
rlabel metal1 1890 1695 1894 1699 1 Add_SubB3
rlabel metal1 3115 1640 3118 1643 1 n3
rlabel metal1 2953 1674 3043 1678 5 VDD
rlabel metal1 3093 1662 3118 1665 1 VDD
rlabel metal1 3093 1625 3118 1628 1 GND
rlabel metal1 2954 1592 3096 1595 1 GND
rlabel metal1 3202 1674 3292 1678 5 VDD
rlabel metal1 3364 1640 3367 1643 1 n2
rlabel metal1 3342 1625 3367 1628 1 GND
rlabel metal1 3342 1662 3367 1665 1 VDD
rlabel metal1 3203 1592 3345 1595 1 GND
rlabel metal1 3459 1674 3549 1678 5 VDD
rlabel metal1 3621 1640 3624 1643 7 n1
rlabel metal1 3599 1662 3624 1665 1 VDD
rlabel metal1 3599 1625 3624 1628 1 GND
rlabel metal1 3460 1592 3602 1595 1 GND
rlabel metal1 3843 1640 3846 1643 7 n0
rlabel metal1 3681 1674 3771 1678 5 VDD
rlabel metal1 3821 1662 3846 1665 1 VDD
rlabel metal1 3821 1625 3846 1628 1 GND
rlabel metal1 3078 1267 3103 1270 1 GND
rlabel metal1 3078 1304 3103 1307 5 VDD
rlabel metal1 3134 1267 3159 1270 1 GND
rlabel metal1 3134 1304 3159 1307 5 VDD
rlabel metal1 3331 1267 3356 1270 1 GND
rlabel metal1 3331 1304 3356 1307 5 VDD
rlabel metal1 3594 1267 3619 1270 1 GND
rlabel metal1 3594 1304 3619 1307 5 VDD
rlabel metal1 3948 1802 4033 1806 5 VDD
rlabel metal1 3943 1769 3947 1773 1 n3
rlabel metal1 3943 1762 3947 1766 1 n2
rlabel metal1 3943 1755 3947 1759 1 n1
rlabel metal1 3943 1748 3947 1752 1 n0
rlabel metal1 4032 1769 4036 1773 1 AEB
rlabel metal1 3997 1426 4074 1430 5 VDD
rlabel metal1 3996 1347 4074 1351 1 GND
rlabel metal1 3994 1395 3998 1399 1 y3
rlabel metal1 3994 1388 3998 1392 1 y2
rlabel metal1 3994 1381 3998 1385 1 y1
rlabel metal1 3994 1374 3998 1378 1 y0
rlabel metal1 4075 1390 4079 1394 7 AGB
rlabel metal1 4279 1608 4283 1612 7 ALB
rlabel metal1 4244 1613 4248 1617 1 AEB
rlabel metal1 4244 1606 4248 1610 1 AGB
rlabel metal1 4247 1644 4281 1649 1 VDD
rlabel metal1 3832 1467 3837 1471 7 y0
rlabel metal1 3731 1467 3736 1471 1 n3
rlabel metal1 3731 1460 3736 1464 1 n2
rlabel metal1 3731 1453 3736 1457 1 n1
rlabel metal1 3294 1448 3299 1452 7 y2
rlabel metal1 3215 1448 3220 1452 1 n3
rlabel metal1 3219 1416 3298 1420 1 GND
rlabel metal1 3220 1481 3297 1485 5 VDD
rlabel metal1 3085 1443 3089 1447 7 y3
rlabel metal1 3017 1415 3086 1418 1 GND
rlabel metal1 3018 1476 3085 1479 5 VDD
rlabel metal1 3475 1490 3560 1493 1 VDD
rlabel metal1 3560 1457 3564 1461 7 y1
rlabel metal1 3470 1450 3474 1454 1 n2
rlabel metal1 3470 1457 3474 1461 1 n3
rlabel metal1 3474 1417 3561 1421 1 GND
rlabel metal1 3013 1443 3017 1447 1 CompA3
rlabel metal1 3013 1434 3017 1438 1 CompB3not
rlabel metal1 3215 1441 3220 1445 1 CompB2not
rlabel metal1 3215 1434 3220 1438 1 CompA2
rlabel metal1 3470 1436 3474 1440 1 CompA1
rlabel metal1 3470 1443 3474 1447 1 CompB1not
rlabel metal1 3731 1438 3736 1442 1 CompB0not
rlabel metal1 3731 1446 3736 1450 1 CompA0
rlabel metal1 3723 1500 3820 1504 1 VDD
rlabel metal1 2947 1632 2951 1636 1 CompA3
rlabel metal1 2948 1624 2952 1628 1 CompB3
rlabel metal1 3194 1624 3198 1628 1 CompB2
rlabel metal1 3194 1632 3198 1636 1 CompA2
rlabel metal1 3451 1632 3455 1636 1 CompA1
rlabel metal1 3451 1624 3455 1628 1 CompB1
rlabel metal1 3673 1632 3677 1636 1 CompA0
rlabel metal1 3678 1624 3680 1628 1 CompB0
rlabel metal1 3078 1282 3081 1286 1 CompB3
rlabel metal1 3095 1282 3098 1285 1 CompB3not
rlabel metal1 3133 1282 3137 1286 1 CompB2
rlabel metal1 3156 1282 3159 1285 1 CompB2not
rlabel metal1 3330 1282 3334 1286 1 CompB1
rlabel metal1 3353 1282 3356 1285 1 CompB1not
rlabel metal1 3593 1282 3597 1286 1 CompB0
rlabel metal1 3616 1282 3619 1285 1 CompB0not
rlabel metal1 3962 1730 3979 1733 1 GND
rlabel space 4319 1705 4326 1718 1 VDD
rlabel space 4390 1671 4397 1684 1 GND
<< end >>
