magic
tech scmos
timestamp 1701512702
<< nwell >>
rect 344 211 434 229
rect 506 220 596 238
rect 743 230 833 248
rect 632 104 669 122
rect 675 104 699 122
rect 760 105 797 123
rect 803 105 827 123
rect 801 33 858 51
rect 353 -121 443 -103
rect 515 -112 605 -94
rect 752 -102 842 -84
rect 641 -228 678 -210
rect 684 -228 708 -210
rect 769 -227 806 -209
rect 812 -227 836 -209
rect 810 -299 867 -281
rect 374 -487 464 -469
rect 536 -478 626 -460
rect 773 -468 863 -450
rect 662 -594 699 -576
rect 705 -594 729 -576
rect 790 -593 827 -575
rect 833 -593 857 -575
rect 831 -665 888 -647
rect 402 -861 492 -843
rect 564 -852 654 -834
rect 801 -842 891 -824
rect 690 -968 727 -950
rect 733 -968 757 -950
rect 818 -967 855 -949
rect 861 -967 885 -949
rect 859 -1039 916 -1021
<< ntransistor >>
rect 355 171 357 175
rect 371 171 373 175
rect 381 171 383 175
rect 391 171 393 175
rect 401 171 403 175
rect 517 180 519 184
rect 533 180 535 184
rect 543 180 545 184
rect 553 180 555 184
rect 563 180 565 184
rect 421 171 423 175
rect 754 190 756 194
rect 770 190 772 194
rect 780 190 782 194
rect 790 190 792 194
rect 800 190 802 194
rect 583 180 585 184
rect 820 190 822 194
rect 643 80 645 84
rect 653 80 655 84
rect 686 80 688 84
rect 771 81 773 85
rect 781 81 783 85
rect 814 81 816 85
rect 812 3 814 7
rect 822 3 824 7
rect 840 3 842 7
rect 364 -161 366 -157
rect 380 -161 382 -157
rect 390 -161 392 -157
rect 400 -161 402 -157
rect 410 -161 412 -157
rect 526 -152 528 -148
rect 542 -152 544 -148
rect 552 -152 554 -148
rect 562 -152 564 -148
rect 572 -152 574 -148
rect 430 -161 432 -157
rect 763 -142 765 -138
rect 779 -142 781 -138
rect 789 -142 791 -138
rect 799 -142 801 -138
rect 809 -142 811 -138
rect 592 -152 594 -148
rect 829 -142 831 -138
rect 652 -252 654 -248
rect 662 -252 664 -248
rect 695 -252 697 -248
rect 780 -251 782 -247
rect 790 -251 792 -247
rect 823 -251 825 -247
rect 821 -329 823 -325
rect 831 -329 833 -325
rect 849 -329 851 -325
rect 385 -527 387 -523
rect 401 -527 403 -523
rect 411 -527 413 -523
rect 421 -527 423 -523
rect 431 -527 433 -523
rect 547 -518 549 -514
rect 563 -518 565 -514
rect 573 -518 575 -514
rect 583 -518 585 -514
rect 593 -518 595 -514
rect 451 -527 453 -523
rect 784 -508 786 -504
rect 800 -508 802 -504
rect 810 -508 812 -504
rect 820 -508 822 -504
rect 830 -508 832 -504
rect 613 -518 615 -514
rect 850 -508 852 -504
rect 673 -618 675 -614
rect 683 -618 685 -614
rect 716 -618 718 -614
rect 801 -617 803 -613
rect 811 -617 813 -613
rect 844 -617 846 -613
rect 842 -695 844 -691
rect 852 -695 854 -691
rect 870 -695 872 -691
rect 413 -901 415 -897
rect 429 -901 431 -897
rect 439 -901 441 -897
rect 449 -901 451 -897
rect 459 -901 461 -897
rect 575 -892 577 -888
rect 591 -892 593 -888
rect 601 -892 603 -888
rect 611 -892 613 -888
rect 621 -892 623 -888
rect 479 -901 481 -897
rect 812 -882 814 -878
rect 828 -882 830 -878
rect 838 -882 840 -878
rect 848 -882 850 -878
rect 858 -882 860 -878
rect 641 -892 643 -888
rect 878 -882 880 -878
rect 701 -992 703 -988
rect 711 -992 713 -988
rect 744 -992 746 -988
rect 829 -991 831 -987
rect 839 -991 841 -987
rect 872 -991 874 -987
rect 870 -1069 872 -1065
rect 880 -1069 882 -1065
rect 898 -1069 900 -1065
<< ptransistor >>
rect 355 217 357 223
rect 371 217 373 223
rect 381 217 383 223
rect 391 217 393 223
rect 401 217 403 223
rect 421 217 423 223
rect 517 226 519 232
rect 533 226 535 232
rect 543 226 545 232
rect 553 226 555 232
rect 563 226 565 232
rect 583 226 585 232
rect 754 236 756 242
rect 770 236 772 242
rect 780 236 782 242
rect 790 236 792 242
rect 800 236 802 242
rect 820 236 822 242
rect 643 110 645 116
rect 653 110 655 116
rect 686 110 688 116
rect 771 111 773 117
rect 781 111 783 117
rect 814 111 816 117
rect 812 39 814 45
rect 822 39 824 45
rect 840 39 842 45
rect 364 -115 366 -109
rect 380 -115 382 -109
rect 390 -115 392 -109
rect 400 -115 402 -109
rect 410 -115 412 -109
rect 430 -115 432 -109
rect 526 -106 528 -100
rect 542 -106 544 -100
rect 552 -106 554 -100
rect 562 -106 564 -100
rect 572 -106 574 -100
rect 592 -106 594 -100
rect 763 -96 765 -90
rect 779 -96 781 -90
rect 789 -96 791 -90
rect 799 -96 801 -90
rect 809 -96 811 -90
rect 829 -96 831 -90
rect 652 -222 654 -216
rect 662 -222 664 -216
rect 695 -222 697 -216
rect 780 -221 782 -215
rect 790 -221 792 -215
rect 823 -221 825 -215
rect 821 -293 823 -287
rect 831 -293 833 -287
rect 849 -293 851 -287
rect 385 -481 387 -475
rect 401 -481 403 -475
rect 411 -481 413 -475
rect 421 -481 423 -475
rect 431 -481 433 -475
rect 451 -481 453 -475
rect 547 -472 549 -466
rect 563 -472 565 -466
rect 573 -472 575 -466
rect 583 -472 585 -466
rect 593 -472 595 -466
rect 613 -472 615 -466
rect 784 -462 786 -456
rect 800 -462 802 -456
rect 810 -462 812 -456
rect 820 -462 822 -456
rect 830 -462 832 -456
rect 850 -462 852 -456
rect 673 -588 675 -582
rect 683 -588 685 -582
rect 716 -588 718 -582
rect 801 -587 803 -581
rect 811 -587 813 -581
rect 844 -587 846 -581
rect 842 -659 844 -653
rect 852 -659 854 -653
rect 870 -659 872 -653
rect 413 -855 415 -849
rect 429 -855 431 -849
rect 439 -855 441 -849
rect 449 -855 451 -849
rect 459 -855 461 -849
rect 479 -855 481 -849
rect 575 -846 577 -840
rect 591 -846 593 -840
rect 601 -846 603 -840
rect 611 -846 613 -840
rect 621 -846 623 -840
rect 641 -846 643 -840
rect 812 -836 814 -830
rect 828 -836 830 -830
rect 838 -836 840 -830
rect 848 -836 850 -830
rect 858 -836 860 -830
rect 878 -836 880 -830
rect 701 -962 703 -956
rect 711 -962 713 -956
rect 744 -962 746 -956
rect 829 -961 831 -955
rect 839 -961 841 -955
rect 872 -961 874 -955
rect 870 -1033 872 -1027
rect 880 -1033 882 -1027
rect 898 -1033 900 -1027
<< ndiffusion >>
rect 354 171 355 175
rect 357 171 358 175
rect 370 171 371 175
rect 373 171 381 175
rect 383 171 385 175
rect 389 171 391 175
rect 393 171 401 175
rect 403 171 404 175
rect 516 180 517 184
rect 519 180 520 184
rect 532 180 533 184
rect 535 180 543 184
rect 545 180 547 184
rect 551 180 553 184
rect 555 180 563 184
rect 565 180 566 184
rect 420 171 421 175
rect 423 171 424 175
rect 753 190 754 194
rect 756 190 757 194
rect 769 190 770 194
rect 772 190 780 194
rect 782 190 784 194
rect 788 190 790 194
rect 792 190 800 194
rect 802 190 803 194
rect 582 180 583 184
rect 585 180 586 184
rect 819 190 820 194
rect 822 190 823 194
rect 642 80 643 84
rect 645 80 653 84
rect 655 80 657 84
rect 685 80 686 84
rect 688 80 689 84
rect 770 81 771 85
rect 773 81 781 85
rect 783 81 785 85
rect 813 81 814 85
rect 816 81 817 85
rect 811 3 812 7
rect 814 3 816 7
rect 820 3 822 7
rect 824 3 825 7
rect 839 3 840 7
rect 842 3 843 7
rect 363 -161 364 -157
rect 366 -161 367 -157
rect 379 -161 380 -157
rect 382 -161 390 -157
rect 392 -161 394 -157
rect 398 -161 400 -157
rect 402 -161 410 -157
rect 412 -161 413 -157
rect 525 -152 526 -148
rect 528 -152 529 -148
rect 541 -152 542 -148
rect 544 -152 552 -148
rect 554 -152 556 -148
rect 560 -152 562 -148
rect 564 -152 572 -148
rect 574 -152 575 -148
rect 429 -161 430 -157
rect 432 -161 433 -157
rect 762 -142 763 -138
rect 765 -142 766 -138
rect 778 -142 779 -138
rect 781 -142 789 -138
rect 791 -142 793 -138
rect 797 -142 799 -138
rect 801 -142 809 -138
rect 811 -142 812 -138
rect 591 -152 592 -148
rect 594 -152 595 -148
rect 828 -142 829 -138
rect 831 -142 832 -138
rect 651 -252 652 -248
rect 654 -252 662 -248
rect 664 -252 666 -248
rect 694 -252 695 -248
rect 697 -252 698 -248
rect 779 -251 780 -247
rect 782 -251 790 -247
rect 792 -251 794 -247
rect 822 -251 823 -247
rect 825 -251 826 -247
rect 820 -329 821 -325
rect 823 -329 825 -325
rect 829 -329 831 -325
rect 833 -329 834 -325
rect 848 -329 849 -325
rect 851 -329 852 -325
rect 384 -527 385 -523
rect 387 -527 388 -523
rect 400 -527 401 -523
rect 403 -527 411 -523
rect 413 -527 415 -523
rect 419 -527 421 -523
rect 423 -527 431 -523
rect 433 -527 434 -523
rect 546 -518 547 -514
rect 549 -518 550 -514
rect 562 -518 563 -514
rect 565 -518 573 -514
rect 575 -518 577 -514
rect 581 -518 583 -514
rect 585 -518 593 -514
rect 595 -518 596 -514
rect 450 -527 451 -523
rect 453 -527 454 -523
rect 783 -508 784 -504
rect 786 -508 787 -504
rect 799 -508 800 -504
rect 802 -508 810 -504
rect 812 -508 814 -504
rect 818 -508 820 -504
rect 822 -508 830 -504
rect 832 -508 833 -504
rect 612 -518 613 -514
rect 615 -518 616 -514
rect 849 -508 850 -504
rect 852 -508 853 -504
rect 672 -618 673 -614
rect 675 -618 683 -614
rect 685 -618 687 -614
rect 715 -618 716 -614
rect 718 -618 719 -614
rect 800 -617 801 -613
rect 803 -617 811 -613
rect 813 -617 815 -613
rect 843 -617 844 -613
rect 846 -617 847 -613
rect 841 -695 842 -691
rect 844 -695 846 -691
rect 850 -695 852 -691
rect 854 -695 855 -691
rect 869 -695 870 -691
rect 872 -695 873 -691
rect 412 -901 413 -897
rect 415 -901 416 -897
rect 428 -901 429 -897
rect 431 -901 439 -897
rect 441 -901 443 -897
rect 447 -901 449 -897
rect 451 -901 459 -897
rect 461 -901 462 -897
rect 574 -892 575 -888
rect 577 -892 578 -888
rect 590 -892 591 -888
rect 593 -892 601 -888
rect 603 -892 605 -888
rect 609 -892 611 -888
rect 613 -892 621 -888
rect 623 -892 624 -888
rect 478 -901 479 -897
rect 481 -901 482 -897
rect 811 -882 812 -878
rect 814 -882 815 -878
rect 827 -882 828 -878
rect 830 -882 838 -878
rect 840 -882 842 -878
rect 846 -882 848 -878
rect 850 -882 858 -878
rect 860 -882 861 -878
rect 640 -892 641 -888
rect 643 -892 644 -888
rect 877 -882 878 -878
rect 880 -882 881 -878
rect 700 -992 701 -988
rect 703 -992 711 -988
rect 713 -992 715 -988
rect 743 -992 744 -988
rect 746 -992 747 -988
rect 828 -991 829 -987
rect 831 -991 839 -987
rect 841 -991 843 -987
rect 871 -991 872 -987
rect 874 -991 875 -987
rect 869 -1069 870 -1065
rect 872 -1069 874 -1065
rect 878 -1069 880 -1065
rect 882 -1069 883 -1065
rect 897 -1069 898 -1065
rect 900 -1069 901 -1065
<< pdiffusion >>
rect 354 217 355 223
rect 357 217 358 223
rect 370 217 371 223
rect 373 217 381 223
rect 383 217 385 223
rect 389 217 391 223
rect 393 217 401 223
rect 403 217 404 223
rect 420 217 421 223
rect 423 217 424 223
rect 516 226 517 232
rect 519 226 520 232
rect 532 226 533 232
rect 535 226 543 232
rect 545 226 547 232
rect 551 226 553 232
rect 555 226 563 232
rect 565 226 566 232
rect 582 226 583 232
rect 585 226 586 232
rect 753 236 754 242
rect 756 236 757 242
rect 769 236 770 242
rect 772 236 780 242
rect 782 236 784 242
rect 788 236 790 242
rect 792 236 800 242
rect 802 236 803 242
rect 819 236 820 242
rect 822 236 823 242
rect 642 110 643 116
rect 645 110 647 116
rect 651 110 653 116
rect 655 110 657 116
rect 685 110 686 116
rect 688 110 689 116
rect 770 111 771 117
rect 773 111 775 117
rect 779 111 781 117
rect 783 111 785 117
rect 813 111 814 117
rect 816 111 817 117
rect 811 39 812 45
rect 814 39 822 45
rect 824 39 825 45
rect 839 39 840 45
rect 842 39 843 45
rect 363 -115 364 -109
rect 366 -115 367 -109
rect 379 -115 380 -109
rect 382 -115 390 -109
rect 392 -115 394 -109
rect 398 -115 400 -109
rect 402 -115 410 -109
rect 412 -115 413 -109
rect 429 -115 430 -109
rect 432 -115 433 -109
rect 525 -106 526 -100
rect 528 -106 529 -100
rect 541 -106 542 -100
rect 544 -106 552 -100
rect 554 -106 556 -100
rect 560 -106 562 -100
rect 564 -106 572 -100
rect 574 -106 575 -100
rect 591 -106 592 -100
rect 594 -106 595 -100
rect 762 -96 763 -90
rect 765 -96 766 -90
rect 778 -96 779 -90
rect 781 -96 789 -90
rect 791 -96 793 -90
rect 797 -96 799 -90
rect 801 -96 809 -90
rect 811 -96 812 -90
rect 828 -96 829 -90
rect 831 -96 832 -90
rect 651 -222 652 -216
rect 654 -222 656 -216
rect 660 -222 662 -216
rect 664 -222 666 -216
rect 694 -222 695 -216
rect 697 -222 698 -216
rect 779 -221 780 -215
rect 782 -221 784 -215
rect 788 -221 790 -215
rect 792 -221 794 -215
rect 822 -221 823 -215
rect 825 -221 826 -215
rect 820 -293 821 -287
rect 823 -293 831 -287
rect 833 -293 834 -287
rect 848 -293 849 -287
rect 851 -293 852 -287
rect 384 -481 385 -475
rect 387 -481 388 -475
rect 400 -481 401 -475
rect 403 -481 411 -475
rect 413 -481 415 -475
rect 419 -481 421 -475
rect 423 -481 431 -475
rect 433 -481 434 -475
rect 450 -481 451 -475
rect 453 -481 454 -475
rect 546 -472 547 -466
rect 549 -472 550 -466
rect 562 -472 563 -466
rect 565 -472 573 -466
rect 575 -472 577 -466
rect 581 -472 583 -466
rect 585 -472 593 -466
rect 595 -472 596 -466
rect 612 -472 613 -466
rect 615 -472 616 -466
rect 783 -462 784 -456
rect 786 -462 787 -456
rect 799 -462 800 -456
rect 802 -462 810 -456
rect 812 -462 814 -456
rect 818 -462 820 -456
rect 822 -462 830 -456
rect 832 -462 833 -456
rect 849 -462 850 -456
rect 852 -462 853 -456
rect 672 -588 673 -582
rect 675 -588 677 -582
rect 681 -588 683 -582
rect 685 -588 687 -582
rect 715 -588 716 -582
rect 718 -588 719 -582
rect 800 -587 801 -581
rect 803 -587 805 -581
rect 809 -587 811 -581
rect 813 -587 815 -581
rect 843 -587 844 -581
rect 846 -587 847 -581
rect 841 -659 842 -653
rect 844 -659 852 -653
rect 854 -659 855 -653
rect 869 -659 870 -653
rect 872 -659 873 -653
rect 412 -855 413 -849
rect 415 -855 416 -849
rect 428 -855 429 -849
rect 431 -855 439 -849
rect 441 -855 443 -849
rect 447 -855 449 -849
rect 451 -855 459 -849
rect 461 -855 462 -849
rect 478 -855 479 -849
rect 481 -855 482 -849
rect 574 -846 575 -840
rect 577 -846 578 -840
rect 590 -846 591 -840
rect 593 -846 601 -840
rect 603 -846 605 -840
rect 609 -846 611 -840
rect 613 -846 621 -840
rect 623 -846 624 -840
rect 640 -846 641 -840
rect 643 -846 644 -840
rect 811 -836 812 -830
rect 814 -836 815 -830
rect 827 -836 828 -830
rect 830 -836 838 -830
rect 840 -836 842 -830
rect 846 -836 848 -830
rect 850 -836 858 -830
rect 860 -836 861 -830
rect 877 -836 878 -830
rect 880 -836 881 -830
rect 700 -962 701 -956
rect 703 -962 705 -956
rect 709 -962 711 -956
rect 713 -962 715 -956
rect 743 -962 744 -956
rect 746 -962 747 -956
rect 828 -961 829 -955
rect 831 -961 833 -955
rect 837 -961 839 -955
rect 841 -961 843 -955
rect 871 -961 872 -955
rect 874 -961 875 -955
rect 869 -1033 870 -1027
rect 872 -1033 880 -1027
rect 882 -1033 883 -1027
rect 897 -1033 898 -1027
rect 900 -1033 901 -1027
<< ndcontact >>
rect 350 171 354 175
rect 358 171 362 175
rect 366 171 370 175
rect 385 171 389 175
rect 404 171 408 175
rect 512 180 516 184
rect 520 180 524 184
rect 528 180 532 184
rect 547 180 551 184
rect 566 180 570 184
rect 416 171 420 175
rect 424 171 428 175
rect 749 190 753 194
rect 757 190 761 194
rect 765 190 769 194
rect 784 190 788 194
rect 803 190 807 194
rect 578 180 582 184
rect 586 180 590 184
rect 815 190 819 194
rect 823 190 827 194
rect 638 80 642 84
rect 657 80 661 84
rect 681 80 685 84
rect 689 80 693 84
rect 766 81 770 85
rect 785 81 789 85
rect 809 81 813 85
rect 817 81 821 85
rect 807 3 811 7
rect 816 3 820 7
rect 825 3 829 7
rect 835 3 839 7
rect 843 3 847 7
rect 359 -161 363 -157
rect 367 -161 371 -157
rect 375 -161 379 -157
rect 394 -161 398 -157
rect 413 -161 417 -157
rect 521 -152 525 -148
rect 529 -152 533 -148
rect 537 -152 541 -148
rect 556 -152 560 -148
rect 575 -152 579 -148
rect 425 -161 429 -157
rect 433 -161 437 -157
rect 758 -142 762 -138
rect 766 -142 770 -138
rect 774 -142 778 -138
rect 793 -142 797 -138
rect 812 -142 816 -138
rect 587 -152 591 -148
rect 595 -152 599 -148
rect 824 -142 828 -138
rect 832 -142 836 -138
rect 647 -252 651 -248
rect 666 -252 670 -248
rect 690 -252 694 -248
rect 698 -252 702 -248
rect 775 -251 779 -247
rect 794 -251 798 -247
rect 818 -251 822 -247
rect 826 -251 830 -247
rect 816 -329 820 -325
rect 825 -329 829 -325
rect 834 -329 838 -325
rect 844 -329 848 -325
rect 852 -329 856 -325
rect 380 -527 384 -523
rect 388 -527 392 -523
rect 396 -527 400 -523
rect 415 -527 419 -523
rect 434 -527 438 -523
rect 542 -518 546 -514
rect 550 -518 554 -514
rect 558 -518 562 -514
rect 577 -518 581 -514
rect 596 -518 600 -514
rect 446 -527 450 -523
rect 454 -527 458 -523
rect 779 -508 783 -504
rect 787 -508 791 -504
rect 795 -508 799 -504
rect 814 -508 818 -504
rect 833 -508 837 -504
rect 608 -518 612 -514
rect 616 -518 620 -514
rect 845 -508 849 -504
rect 853 -508 857 -504
rect 668 -618 672 -614
rect 687 -618 691 -614
rect 711 -618 715 -614
rect 719 -618 723 -614
rect 796 -617 800 -613
rect 815 -617 819 -613
rect 839 -617 843 -613
rect 847 -617 851 -613
rect 837 -695 841 -691
rect 846 -695 850 -691
rect 855 -695 859 -691
rect 865 -695 869 -691
rect 873 -695 877 -691
rect 408 -901 412 -897
rect 416 -901 420 -897
rect 424 -901 428 -897
rect 443 -901 447 -897
rect 462 -901 466 -897
rect 570 -892 574 -888
rect 578 -892 582 -888
rect 586 -892 590 -888
rect 605 -892 609 -888
rect 624 -892 628 -888
rect 474 -901 478 -897
rect 482 -901 486 -897
rect 807 -882 811 -878
rect 815 -882 819 -878
rect 823 -882 827 -878
rect 842 -882 846 -878
rect 861 -882 865 -878
rect 636 -892 640 -888
rect 644 -892 648 -888
rect 873 -882 877 -878
rect 881 -882 885 -878
rect 696 -992 700 -988
rect 715 -992 719 -988
rect 739 -992 743 -988
rect 747 -992 751 -988
rect 824 -991 828 -987
rect 843 -991 847 -987
rect 867 -991 871 -987
rect 875 -991 879 -987
rect 865 -1069 869 -1065
rect 874 -1069 878 -1065
rect 883 -1069 887 -1065
rect 893 -1069 897 -1065
rect 901 -1069 905 -1065
<< pdcontact >>
rect 350 217 354 223
rect 358 217 362 223
rect 366 217 370 223
rect 385 217 389 223
rect 404 217 408 223
rect 416 217 420 223
rect 424 217 428 223
rect 512 226 516 232
rect 520 226 524 232
rect 528 226 532 232
rect 547 226 551 232
rect 566 226 570 232
rect 578 226 582 232
rect 586 226 590 232
rect 749 236 753 242
rect 757 236 761 242
rect 765 236 769 242
rect 784 236 788 242
rect 803 236 807 242
rect 815 236 819 242
rect 823 236 827 242
rect 638 110 642 116
rect 647 110 651 116
rect 657 110 661 116
rect 681 110 685 116
rect 689 110 693 116
rect 766 111 770 117
rect 775 111 779 117
rect 785 111 789 117
rect 809 111 813 117
rect 817 111 821 117
rect 807 39 811 45
rect 825 39 829 45
rect 835 39 839 45
rect 843 39 847 45
rect 359 -115 363 -109
rect 367 -115 371 -109
rect 375 -115 379 -109
rect 394 -115 398 -109
rect 413 -115 417 -109
rect 425 -115 429 -109
rect 433 -115 437 -109
rect 521 -106 525 -100
rect 529 -106 533 -100
rect 537 -106 541 -100
rect 556 -106 560 -100
rect 575 -106 579 -100
rect 587 -106 591 -100
rect 595 -106 599 -100
rect 758 -96 762 -90
rect 766 -96 770 -90
rect 774 -96 778 -90
rect 793 -96 797 -90
rect 812 -96 816 -90
rect 824 -96 828 -90
rect 832 -96 836 -90
rect 647 -222 651 -216
rect 656 -222 660 -216
rect 666 -222 670 -216
rect 690 -222 694 -216
rect 698 -222 702 -216
rect 775 -221 779 -215
rect 784 -221 788 -215
rect 794 -221 798 -215
rect 818 -221 822 -215
rect 826 -221 830 -215
rect 816 -293 820 -287
rect 834 -293 838 -287
rect 844 -293 848 -287
rect 852 -293 856 -287
rect 380 -481 384 -475
rect 388 -481 392 -475
rect 396 -481 400 -475
rect 415 -481 419 -475
rect 434 -481 438 -475
rect 446 -481 450 -475
rect 454 -481 458 -475
rect 542 -472 546 -466
rect 550 -472 554 -466
rect 558 -472 562 -466
rect 577 -472 581 -466
rect 596 -472 600 -466
rect 608 -472 612 -466
rect 616 -472 620 -466
rect 779 -462 783 -456
rect 787 -462 791 -456
rect 795 -462 799 -456
rect 814 -462 818 -456
rect 833 -462 837 -456
rect 845 -462 849 -456
rect 853 -462 857 -456
rect 668 -588 672 -582
rect 677 -588 681 -582
rect 687 -588 691 -582
rect 711 -588 715 -582
rect 719 -588 723 -582
rect 796 -587 800 -581
rect 805 -587 809 -581
rect 815 -587 819 -581
rect 839 -587 843 -581
rect 847 -587 851 -581
rect 837 -659 841 -653
rect 855 -659 859 -653
rect 865 -659 869 -653
rect 873 -659 877 -653
rect 408 -855 412 -849
rect 416 -855 420 -849
rect 424 -855 428 -849
rect 443 -855 447 -849
rect 462 -855 466 -849
rect 474 -855 478 -849
rect 482 -855 486 -849
rect 570 -846 574 -840
rect 578 -846 582 -840
rect 586 -846 590 -840
rect 605 -846 609 -840
rect 624 -846 628 -840
rect 636 -846 640 -840
rect 644 -846 648 -840
rect 807 -836 811 -830
rect 815 -836 819 -830
rect 823 -836 827 -830
rect 842 -836 846 -830
rect 861 -836 865 -830
rect 873 -836 877 -830
rect 881 -836 885 -830
rect 696 -962 700 -956
rect 705 -962 709 -956
rect 715 -962 719 -956
rect 739 -962 743 -956
rect 747 -962 751 -956
rect 824 -961 828 -955
rect 833 -961 837 -955
rect 843 -961 847 -955
rect 867 -961 871 -955
rect 875 -961 879 -955
rect 865 -1033 869 -1027
rect 883 -1033 887 -1027
rect 893 -1033 897 -1027
rect 901 -1033 905 -1027
<< polysilicon >>
rect 754 250 840 252
rect 754 242 756 250
rect 770 242 772 245
rect 780 242 782 245
rect 790 242 792 250
rect 800 242 802 245
rect 820 242 822 245
rect 517 240 603 242
rect 355 231 441 233
rect 517 232 519 240
rect 533 232 535 235
rect 543 232 545 235
rect 553 232 555 240
rect 563 232 565 235
rect 583 232 585 235
rect 355 223 357 231
rect 371 223 373 226
rect 381 223 383 226
rect 391 223 393 231
rect 401 223 403 226
rect 421 223 423 226
rect 355 175 357 217
rect 371 175 373 217
rect 381 196 383 217
rect 391 214 393 217
rect 381 194 393 196
rect 381 175 383 178
rect 391 175 393 194
rect 401 175 403 217
rect 421 194 423 217
rect 439 189 441 231
rect 412 187 441 189
rect 355 168 357 171
rect 371 160 373 171
rect 381 165 383 171
rect 391 168 393 171
rect 401 168 403 171
rect 412 165 414 187
rect 517 184 519 226
rect 533 184 535 226
rect 543 205 545 226
rect 553 223 555 226
rect 543 203 555 205
rect 543 184 545 187
rect 553 184 555 203
rect 563 184 565 226
rect 583 203 585 226
rect 601 198 603 240
rect 574 196 603 198
rect 421 175 423 183
rect 517 177 519 180
rect 381 163 414 165
rect 421 160 423 171
rect 533 169 535 180
rect 543 174 545 180
rect 553 177 555 180
rect 563 177 565 180
rect 574 174 576 196
rect 754 194 756 236
rect 770 194 772 236
rect 780 215 782 236
rect 790 233 792 236
rect 780 213 792 215
rect 780 194 782 197
rect 790 194 792 213
rect 800 194 802 236
rect 820 213 822 236
rect 838 208 840 250
rect 811 206 840 208
rect 583 184 585 192
rect 754 187 756 190
rect 543 172 576 174
rect 583 169 585 180
rect 770 179 772 190
rect 780 184 782 190
rect 790 187 792 190
rect 800 187 802 190
rect 811 184 813 206
rect 820 194 822 202
rect 780 182 813 184
rect 820 179 822 190
rect 770 177 822 179
rect 533 167 585 169
rect 371 158 423 160
rect 643 116 645 125
rect 653 116 655 125
rect 686 116 688 125
rect 771 117 773 126
rect 781 117 783 126
rect 814 117 816 126
rect 643 84 645 110
rect 653 84 655 110
rect 686 84 688 110
rect 771 85 773 111
rect 781 85 783 111
rect 814 85 816 111
rect 643 77 645 80
rect 653 77 655 80
rect 686 77 688 80
rect 771 78 773 81
rect 781 78 783 81
rect 814 78 816 81
rect 812 45 814 48
rect 822 45 824 48
rect 840 45 842 48
rect 812 7 814 39
rect 822 7 824 39
rect 840 7 842 39
rect 812 0 814 3
rect 822 0 824 3
rect 840 0 842 3
rect 763 -82 849 -80
rect 763 -90 765 -82
rect 779 -90 781 -87
rect 789 -90 791 -87
rect 799 -90 801 -82
rect 809 -90 811 -87
rect 829 -90 831 -87
rect 526 -92 612 -90
rect 364 -101 450 -99
rect 526 -100 528 -92
rect 542 -100 544 -97
rect 552 -100 554 -97
rect 562 -100 564 -92
rect 572 -100 574 -97
rect 592 -100 594 -97
rect 364 -109 366 -101
rect 380 -109 382 -106
rect 390 -109 392 -106
rect 400 -109 402 -101
rect 410 -109 412 -106
rect 430 -109 432 -106
rect 364 -157 366 -115
rect 380 -157 382 -115
rect 390 -136 392 -115
rect 400 -118 402 -115
rect 390 -138 402 -136
rect 390 -157 392 -154
rect 400 -157 402 -138
rect 410 -157 412 -115
rect 430 -138 432 -115
rect 448 -143 450 -101
rect 421 -145 450 -143
rect 364 -164 366 -161
rect 380 -172 382 -161
rect 390 -167 392 -161
rect 400 -164 402 -161
rect 410 -164 412 -161
rect 421 -167 423 -145
rect 526 -148 528 -106
rect 542 -148 544 -106
rect 552 -127 554 -106
rect 562 -109 564 -106
rect 552 -129 564 -127
rect 552 -148 554 -145
rect 562 -148 564 -129
rect 572 -148 574 -106
rect 592 -129 594 -106
rect 610 -134 612 -92
rect 583 -136 612 -134
rect 430 -157 432 -149
rect 526 -155 528 -152
rect 390 -169 423 -167
rect 430 -172 432 -161
rect 542 -163 544 -152
rect 552 -158 554 -152
rect 562 -155 564 -152
rect 572 -155 574 -152
rect 583 -158 585 -136
rect 763 -138 765 -96
rect 779 -138 781 -96
rect 789 -117 791 -96
rect 799 -99 801 -96
rect 789 -119 801 -117
rect 789 -138 791 -135
rect 799 -138 801 -119
rect 809 -138 811 -96
rect 829 -119 831 -96
rect 847 -124 849 -82
rect 820 -126 849 -124
rect 592 -148 594 -140
rect 763 -145 765 -142
rect 552 -160 585 -158
rect 592 -163 594 -152
rect 779 -153 781 -142
rect 789 -148 791 -142
rect 799 -145 801 -142
rect 809 -145 811 -142
rect 820 -148 822 -126
rect 829 -138 831 -130
rect 789 -150 822 -148
rect 829 -153 831 -142
rect 779 -155 831 -153
rect 542 -165 594 -163
rect 380 -174 432 -172
rect 652 -216 654 -207
rect 662 -216 664 -207
rect 695 -216 697 -207
rect 780 -215 782 -206
rect 790 -215 792 -206
rect 823 -215 825 -206
rect 652 -248 654 -222
rect 662 -248 664 -222
rect 695 -248 697 -222
rect 780 -247 782 -221
rect 790 -247 792 -221
rect 823 -247 825 -221
rect 652 -255 654 -252
rect 662 -255 664 -252
rect 695 -255 697 -252
rect 780 -254 782 -251
rect 790 -254 792 -251
rect 823 -254 825 -251
rect 821 -287 823 -284
rect 831 -287 833 -284
rect 849 -287 851 -284
rect 821 -325 823 -293
rect 831 -325 833 -293
rect 849 -325 851 -293
rect 821 -332 823 -329
rect 831 -332 833 -329
rect 849 -332 851 -329
rect 784 -448 870 -446
rect 784 -456 786 -448
rect 800 -456 802 -453
rect 810 -456 812 -453
rect 820 -456 822 -448
rect 830 -456 832 -453
rect 850 -456 852 -453
rect 547 -458 633 -456
rect 385 -467 471 -465
rect 547 -466 549 -458
rect 563 -466 565 -463
rect 573 -466 575 -463
rect 583 -466 585 -458
rect 593 -466 595 -463
rect 613 -466 615 -463
rect 385 -475 387 -467
rect 401 -475 403 -472
rect 411 -475 413 -472
rect 421 -475 423 -467
rect 431 -475 433 -472
rect 451 -475 453 -472
rect 385 -523 387 -481
rect 401 -523 403 -481
rect 411 -502 413 -481
rect 421 -484 423 -481
rect 411 -504 423 -502
rect 411 -523 413 -520
rect 421 -523 423 -504
rect 431 -523 433 -481
rect 451 -504 453 -481
rect 469 -509 471 -467
rect 442 -511 471 -509
rect 385 -530 387 -527
rect 401 -538 403 -527
rect 411 -533 413 -527
rect 421 -530 423 -527
rect 431 -530 433 -527
rect 442 -533 444 -511
rect 547 -514 549 -472
rect 563 -514 565 -472
rect 573 -493 575 -472
rect 583 -475 585 -472
rect 573 -495 585 -493
rect 573 -514 575 -511
rect 583 -514 585 -495
rect 593 -514 595 -472
rect 613 -495 615 -472
rect 631 -500 633 -458
rect 604 -502 633 -500
rect 451 -523 453 -515
rect 547 -521 549 -518
rect 411 -535 444 -533
rect 451 -538 453 -527
rect 563 -529 565 -518
rect 573 -524 575 -518
rect 583 -521 585 -518
rect 593 -521 595 -518
rect 604 -524 606 -502
rect 784 -504 786 -462
rect 800 -504 802 -462
rect 810 -483 812 -462
rect 820 -465 822 -462
rect 810 -485 822 -483
rect 810 -504 812 -501
rect 820 -504 822 -485
rect 830 -504 832 -462
rect 850 -485 852 -462
rect 868 -490 870 -448
rect 841 -492 870 -490
rect 613 -514 615 -506
rect 784 -511 786 -508
rect 573 -526 606 -524
rect 613 -529 615 -518
rect 800 -519 802 -508
rect 810 -514 812 -508
rect 820 -511 822 -508
rect 830 -511 832 -508
rect 841 -514 843 -492
rect 850 -504 852 -496
rect 810 -516 843 -514
rect 850 -519 852 -508
rect 800 -521 852 -519
rect 563 -531 615 -529
rect 401 -540 453 -538
rect 673 -582 675 -573
rect 683 -582 685 -573
rect 716 -582 718 -573
rect 801 -581 803 -572
rect 811 -581 813 -572
rect 844 -581 846 -572
rect 673 -614 675 -588
rect 683 -614 685 -588
rect 716 -614 718 -588
rect 801 -613 803 -587
rect 811 -613 813 -587
rect 844 -613 846 -587
rect 673 -621 675 -618
rect 683 -621 685 -618
rect 716 -621 718 -618
rect 801 -620 803 -617
rect 811 -620 813 -617
rect 844 -620 846 -617
rect 842 -653 844 -650
rect 852 -653 854 -650
rect 870 -653 872 -650
rect 842 -691 844 -659
rect 852 -691 854 -659
rect 870 -691 872 -659
rect 842 -698 844 -695
rect 852 -698 854 -695
rect 870 -698 872 -695
rect 812 -822 898 -820
rect 812 -830 814 -822
rect 828 -830 830 -827
rect 838 -830 840 -827
rect 848 -830 850 -822
rect 858 -830 860 -827
rect 878 -830 880 -827
rect 575 -832 661 -830
rect 413 -841 499 -839
rect 575 -840 577 -832
rect 591 -840 593 -837
rect 601 -840 603 -837
rect 611 -840 613 -832
rect 621 -840 623 -837
rect 641 -840 643 -837
rect 413 -849 415 -841
rect 429 -849 431 -846
rect 439 -849 441 -846
rect 449 -849 451 -841
rect 459 -849 461 -846
rect 479 -849 481 -846
rect 413 -897 415 -855
rect 429 -897 431 -855
rect 439 -876 441 -855
rect 449 -858 451 -855
rect 439 -878 451 -876
rect 439 -897 441 -894
rect 449 -897 451 -878
rect 459 -897 461 -855
rect 479 -878 481 -855
rect 497 -883 499 -841
rect 470 -885 499 -883
rect 413 -904 415 -901
rect 429 -912 431 -901
rect 439 -907 441 -901
rect 449 -904 451 -901
rect 459 -904 461 -901
rect 470 -907 472 -885
rect 575 -888 577 -846
rect 591 -888 593 -846
rect 601 -867 603 -846
rect 611 -849 613 -846
rect 601 -869 613 -867
rect 601 -888 603 -885
rect 611 -888 613 -869
rect 621 -888 623 -846
rect 641 -869 643 -846
rect 659 -874 661 -832
rect 632 -876 661 -874
rect 479 -897 481 -889
rect 575 -895 577 -892
rect 439 -909 472 -907
rect 479 -912 481 -901
rect 591 -903 593 -892
rect 601 -898 603 -892
rect 611 -895 613 -892
rect 621 -895 623 -892
rect 632 -898 634 -876
rect 812 -878 814 -836
rect 828 -878 830 -836
rect 838 -857 840 -836
rect 848 -839 850 -836
rect 838 -859 850 -857
rect 838 -878 840 -875
rect 848 -878 850 -859
rect 858 -878 860 -836
rect 878 -859 880 -836
rect 896 -864 898 -822
rect 869 -866 898 -864
rect 641 -888 643 -880
rect 812 -885 814 -882
rect 601 -900 634 -898
rect 641 -903 643 -892
rect 828 -893 830 -882
rect 838 -888 840 -882
rect 848 -885 850 -882
rect 858 -885 860 -882
rect 869 -888 871 -866
rect 878 -878 880 -870
rect 838 -890 871 -888
rect 878 -893 880 -882
rect 828 -895 880 -893
rect 591 -905 643 -903
rect 429 -914 481 -912
rect 701 -956 703 -947
rect 711 -956 713 -947
rect 744 -956 746 -947
rect 829 -955 831 -946
rect 839 -955 841 -946
rect 872 -955 874 -946
rect 701 -988 703 -962
rect 711 -988 713 -962
rect 744 -988 746 -962
rect 829 -987 831 -961
rect 839 -987 841 -961
rect 872 -987 874 -961
rect 701 -995 703 -992
rect 711 -995 713 -992
rect 744 -995 746 -992
rect 829 -994 831 -991
rect 839 -994 841 -991
rect 872 -994 874 -991
rect 870 -1027 872 -1024
rect 880 -1027 882 -1024
rect 898 -1027 900 -1024
rect 870 -1065 872 -1033
rect 880 -1065 882 -1033
rect 898 -1065 900 -1033
rect 870 -1072 872 -1069
rect 880 -1072 882 -1069
rect 898 -1072 900 -1069
<< polycontact >>
rect 351 194 355 198
rect 377 194 381 198
rect 403 194 407 198
rect 423 194 427 198
rect 513 203 517 207
rect 539 203 543 207
rect 565 203 569 207
rect 585 203 589 207
rect 750 213 754 217
rect 423 179 427 183
rect 776 213 780 217
rect 802 213 806 217
rect 822 213 826 217
rect 585 188 589 192
rect 822 198 826 202
rect 639 98 643 102
rect 649 89 653 93
rect 682 98 686 102
rect 767 99 771 103
rect 777 90 781 94
rect 810 99 814 103
rect 808 26 812 30
rect 818 19 822 23
rect 836 21 840 25
rect 360 -138 364 -134
rect 386 -138 390 -134
rect 412 -138 416 -134
rect 432 -138 436 -134
rect 522 -129 526 -125
rect 548 -129 552 -125
rect 574 -129 578 -125
rect 594 -129 598 -125
rect 759 -119 763 -115
rect 432 -153 436 -149
rect 785 -119 789 -115
rect 811 -119 815 -115
rect 831 -119 835 -115
rect 594 -144 598 -140
rect 831 -134 835 -130
rect 648 -234 652 -230
rect 658 -243 662 -239
rect 691 -234 695 -230
rect 776 -233 780 -229
rect 786 -242 790 -238
rect 819 -233 823 -229
rect 817 -306 821 -302
rect 827 -313 831 -309
rect 845 -311 849 -307
rect 381 -504 385 -500
rect 407 -504 411 -500
rect 433 -504 437 -500
rect 453 -504 457 -500
rect 543 -495 547 -491
rect 569 -495 573 -491
rect 595 -495 599 -491
rect 615 -495 619 -491
rect 780 -485 784 -481
rect 453 -519 457 -515
rect 806 -485 810 -481
rect 832 -485 836 -481
rect 852 -485 856 -481
rect 615 -510 619 -506
rect 852 -500 856 -496
rect 669 -600 673 -596
rect 679 -609 683 -605
rect 712 -600 716 -596
rect 797 -599 801 -595
rect 807 -608 811 -604
rect 840 -599 844 -595
rect 838 -672 842 -668
rect 848 -679 852 -675
rect 866 -677 870 -673
rect 409 -878 413 -874
rect 435 -878 439 -874
rect 461 -878 465 -874
rect 481 -878 485 -874
rect 571 -869 575 -865
rect 597 -869 601 -865
rect 623 -869 627 -865
rect 643 -869 647 -865
rect 808 -859 812 -855
rect 481 -893 485 -889
rect 834 -859 838 -855
rect 860 -859 864 -855
rect 880 -859 884 -855
rect 643 -884 647 -880
rect 880 -874 884 -870
rect 697 -974 701 -970
rect 707 -983 711 -979
rect 740 -974 744 -970
rect 825 -973 829 -969
rect 835 -982 839 -978
rect 868 -973 872 -969
rect 866 -1046 870 -1042
rect 876 -1053 880 -1049
rect 894 -1051 898 -1047
<< metal1 >>
rect 1032 291 1040 292
rect 861 285 1040 291
rect 861 259 866 285
rect 714 255 874 259
rect 714 250 719 255
rect 592 249 719 250
rect 478 245 719 249
rect 478 240 482 245
rect 344 236 482 240
rect 350 223 354 236
rect 366 223 370 236
rect 404 223 408 236
rect 424 223 428 236
rect 512 232 516 245
rect 528 232 532 245
rect 566 232 570 245
rect 586 232 590 245
rect 749 242 753 255
rect 765 242 769 255
rect 803 242 807 255
rect 823 242 827 255
rect 358 198 362 217
rect 385 207 389 217
rect 270 194 351 198
rect 358 194 377 198
rect 270 103 276 194
rect 336 186 344 190
rect 358 175 362 194
rect 385 175 389 202
rect 416 198 420 217
rect 520 207 524 226
rect 547 216 551 226
rect 458 206 513 207
rect 451 203 513 206
rect 520 203 539 207
rect 451 202 487 203
rect 407 194 420 198
rect 416 175 420 194
rect 427 191 431 198
rect 458 193 464 199
rect 427 179 431 186
rect 350 157 354 171
rect 366 157 370 171
rect 404 157 408 171
rect 424 157 428 171
rect 345 153 430 157
rect 458 103 463 157
rect 269 98 464 103
rect 481 102 487 202
rect 499 195 506 199
rect 499 194 503 195
rect 520 184 524 203
rect 547 184 551 211
rect 578 207 582 226
rect 618 215 726 217
rect 613 213 726 215
rect 757 217 761 236
rect 784 226 788 236
rect 731 213 750 217
rect 757 213 776 217
rect 613 211 622 213
rect 569 203 582 207
rect 578 184 582 203
rect 589 200 593 207
rect 589 188 593 195
rect 719 205 743 209
rect 512 166 516 180
rect 528 166 532 180
rect 566 166 570 180
rect 586 166 590 180
rect 598 166 603 168
rect 507 162 603 166
rect 719 156 723 205
rect 757 194 761 213
rect 784 194 788 221
rect 815 217 819 236
rect 896 221 902 226
rect 806 213 819 217
rect 815 194 819 213
rect 826 210 830 217
rect 826 198 830 205
rect 749 176 753 190
rect 765 176 769 190
rect 803 176 807 190
rect 823 176 827 190
rect 749 172 993 176
rect 512 152 723 156
rect 632 131 696 134
rect 638 116 642 131
rect 657 116 661 131
rect 681 116 685 131
rect 647 102 651 110
rect 689 102 693 110
rect 719 103 723 152
rect 763 132 851 135
rect 766 117 770 132
rect 785 117 789 132
rect 809 117 813 132
rect 859 132 874 135
rect 775 103 779 111
rect 817 103 821 111
rect 699 102 712 103
rect 481 98 639 102
rect 647 98 682 102
rect 689 98 712 102
rect 719 99 767 103
rect 775 99 810 103
rect 817 99 874 103
rect 270 -134 276 98
rect 482 97 631 98
rect 611 89 649 93
rect 657 84 661 98
rect 689 84 693 98
rect 608 73 633 74
rect 638 73 642 80
rect 681 73 685 80
rect 608 70 695 73
rect 705 23 712 98
rect 731 90 777 94
rect 785 85 789 99
rect 817 85 821 99
rect 766 74 770 81
rect 809 74 813 81
rect 763 71 828 74
rect 801 57 851 62
rect 807 45 811 57
rect 835 45 839 57
rect 761 26 808 30
rect 761 -18 765 26
rect 825 25 829 39
rect 843 25 847 39
rect 804 19 818 23
rect 825 21 836 25
rect 843 21 859 25
rect 825 15 829 21
rect 816 11 829 15
rect 816 7 820 11
rect 843 7 847 21
rect 807 -4 811 3
rect 825 -4 829 3
rect 835 -4 839 3
rect 803 -9 852 -4
rect 870 -18 874 99
rect 761 -23 874 -18
rect 898 -32 903 26
rect 987 -4 993 172
rect 723 -77 868 -73
rect 873 -77 883 -73
rect 723 -82 728 -77
rect 601 -83 728 -82
rect 493 -87 728 -83
rect 493 -92 497 -87
rect 353 -96 497 -92
rect 359 -109 363 -96
rect 375 -109 379 -96
rect 413 -109 417 -96
rect 433 -109 437 -96
rect 521 -100 525 -87
rect 537 -100 541 -87
rect 575 -100 579 -87
rect 595 -100 599 -87
rect 758 -90 762 -77
rect 774 -90 778 -77
rect 812 -90 816 -77
rect 832 -90 836 -77
rect 367 -134 371 -115
rect 394 -125 398 -115
rect 270 -138 360 -134
rect 367 -138 386 -134
rect 270 -500 276 -138
rect 345 -146 353 -142
rect 367 -157 371 -138
rect 394 -157 398 -130
rect 425 -134 429 -115
rect 529 -125 533 -106
rect 556 -116 560 -106
rect 467 -126 522 -125
rect 460 -129 522 -126
rect 529 -129 548 -125
rect 460 -130 496 -129
rect 416 -138 429 -134
rect 425 -157 429 -138
rect 436 -141 440 -134
rect 467 -139 473 -133
rect 436 -153 440 -146
rect 359 -175 363 -161
rect 375 -175 379 -161
rect 413 -175 417 -161
rect 433 -175 437 -161
rect 354 -179 442 -175
rect 467 -181 472 -175
rect 490 -230 496 -130
rect 508 -137 515 -133
rect 508 -138 512 -137
rect 529 -148 533 -129
rect 556 -148 560 -121
rect 587 -125 591 -106
rect 627 -117 735 -115
rect 622 -119 735 -117
rect 766 -115 770 -96
rect 793 -106 797 -96
rect 740 -119 759 -115
rect 766 -119 785 -115
rect 622 -121 631 -119
rect 578 -129 591 -125
rect 587 -148 591 -129
rect 598 -132 602 -125
rect 598 -144 602 -137
rect 728 -127 752 -123
rect 521 -166 525 -152
rect 537 -166 541 -152
rect 575 -166 579 -152
rect 595 -166 599 -152
rect 607 -166 612 -164
rect 516 -170 612 -166
rect 728 -176 732 -127
rect 766 -138 770 -119
rect 793 -138 797 -111
rect 824 -115 828 -96
rect 905 -111 911 -106
rect 815 -119 828 -115
rect 824 -138 828 -119
rect 835 -122 839 -115
rect 835 -134 839 -127
rect 758 -156 762 -142
rect 774 -156 778 -142
rect 812 -156 816 -142
rect 832 -156 836 -142
rect 758 -160 843 -156
rect 521 -180 732 -176
rect 641 -201 705 -198
rect 647 -216 651 -201
rect 666 -216 670 -201
rect 690 -216 694 -201
rect 656 -230 660 -222
rect 698 -230 702 -222
rect 728 -229 732 -180
rect 772 -200 860 -197
rect 775 -215 779 -200
rect 794 -215 798 -200
rect 818 -215 822 -200
rect 868 -200 883 -197
rect 784 -229 788 -221
rect 826 -229 830 -221
rect 708 -230 721 -229
rect 490 -234 648 -230
rect 656 -234 691 -230
rect 698 -234 721 -230
rect 728 -233 776 -229
rect 784 -233 819 -229
rect 826 -233 883 -229
rect 491 -235 649 -234
rect 620 -243 658 -239
rect 666 -248 670 -234
rect 698 -248 702 -234
rect 617 -259 642 -258
rect 647 -259 651 -252
rect 690 -259 694 -252
rect 617 -262 704 -259
rect 714 -309 721 -234
rect 740 -242 786 -238
rect 794 -247 798 -233
rect 826 -247 830 -233
rect 775 -258 779 -251
rect 818 -258 822 -251
rect 772 -261 837 -258
rect 810 -275 860 -270
rect 816 -287 820 -275
rect 844 -287 848 -275
rect 770 -306 817 -302
rect 770 -350 774 -306
rect 834 -307 838 -293
rect 852 -307 856 -293
rect 813 -313 827 -309
rect 834 -311 845 -307
rect 852 -311 868 -307
rect 834 -317 838 -311
rect 825 -321 838 -317
rect 825 -325 829 -321
rect 852 -325 856 -311
rect 816 -336 820 -329
rect 834 -336 838 -329
rect 844 -336 848 -329
rect 812 -341 866 -336
rect 879 -350 883 -233
rect 770 -355 883 -350
rect 907 -398 912 -306
rect 987 -336 993 -9
rect 1032 -58 1040 285
rect 884 -439 888 -434
rect 744 -443 904 -439
rect 744 -448 749 -443
rect 622 -449 749 -448
rect 516 -453 749 -449
rect 517 -458 521 -453
rect 374 -462 521 -458
rect 380 -475 384 -462
rect 396 -475 400 -462
rect 434 -475 438 -462
rect 454 -475 458 -462
rect 542 -466 546 -453
rect 558 -466 562 -453
rect 596 -466 600 -453
rect 616 -466 620 -453
rect 779 -456 783 -443
rect 795 -456 799 -443
rect 833 -456 837 -443
rect 853 -456 857 -443
rect 388 -500 392 -481
rect 415 -491 419 -481
rect 269 -504 381 -500
rect 388 -504 407 -500
rect 270 -882 276 -504
rect 366 -512 374 -508
rect 388 -523 392 -504
rect 415 -523 419 -496
rect 446 -500 450 -481
rect 550 -491 554 -472
rect 577 -482 581 -472
rect 488 -492 543 -491
rect 481 -495 543 -492
rect 550 -495 569 -491
rect 481 -496 517 -495
rect 437 -504 450 -500
rect 446 -523 450 -504
rect 457 -507 461 -500
rect 488 -505 494 -499
rect 457 -519 461 -512
rect 380 -541 384 -527
rect 396 -541 400 -527
rect 434 -541 438 -527
rect 454 -541 458 -527
rect 375 -545 461 -541
rect 488 -547 493 -541
rect 511 -596 517 -496
rect 529 -503 536 -499
rect 529 -504 533 -503
rect 550 -514 554 -495
rect 577 -514 581 -487
rect 608 -491 612 -472
rect 648 -483 756 -481
rect 643 -485 756 -483
rect 787 -481 791 -462
rect 814 -472 818 -462
rect 761 -485 780 -481
rect 787 -485 806 -481
rect 643 -487 652 -485
rect 599 -495 612 -491
rect 608 -514 612 -495
rect 619 -498 623 -491
rect 619 -510 623 -503
rect 749 -493 773 -489
rect 542 -532 546 -518
rect 558 -532 562 -518
rect 596 -532 600 -518
rect 616 -532 620 -518
rect 628 -532 633 -530
rect 537 -536 633 -532
rect 749 -542 753 -493
rect 787 -504 791 -485
rect 814 -504 818 -477
rect 845 -481 849 -462
rect 926 -477 932 -472
rect 836 -485 849 -481
rect 845 -504 849 -485
rect 856 -488 860 -481
rect 856 -500 860 -493
rect 779 -522 783 -508
rect 795 -522 799 -508
rect 833 -522 837 -508
rect 853 -522 857 -508
rect 779 -526 864 -522
rect 542 -546 753 -542
rect 662 -567 726 -564
rect 668 -582 672 -567
rect 687 -582 691 -567
rect 711 -582 715 -567
rect 677 -596 681 -588
rect 719 -596 723 -588
rect 749 -595 753 -546
rect 793 -566 881 -563
rect 796 -581 800 -566
rect 815 -581 819 -566
rect 839 -581 843 -566
rect 889 -566 904 -563
rect 805 -595 809 -587
rect 847 -595 851 -587
rect 729 -596 742 -595
rect 511 -600 669 -596
rect 677 -600 712 -596
rect 719 -600 742 -596
rect 749 -599 797 -595
rect 805 -599 840 -595
rect 847 -599 904 -595
rect 512 -601 661 -600
rect 641 -609 679 -605
rect 687 -614 691 -600
rect 719 -614 723 -600
rect 638 -625 663 -624
rect 668 -625 672 -618
rect 711 -625 715 -618
rect 638 -628 725 -625
rect 735 -675 742 -600
rect 761 -608 807 -604
rect 815 -613 819 -599
rect 847 -613 851 -599
rect 796 -624 800 -617
rect 839 -624 843 -617
rect 793 -627 858 -624
rect 831 -641 881 -636
rect 837 -653 841 -641
rect 865 -653 869 -641
rect 791 -672 838 -668
rect 791 -716 795 -672
rect 855 -673 859 -659
rect 873 -673 877 -659
rect 834 -679 848 -675
rect 855 -677 866 -673
rect 873 -677 889 -673
rect 855 -683 859 -677
rect 846 -687 859 -683
rect 846 -691 850 -687
rect 873 -691 877 -677
rect 837 -702 841 -695
rect 855 -702 859 -695
rect 865 -702 869 -695
rect 833 -707 887 -702
rect 900 -716 904 -599
rect 791 -721 904 -716
rect 928 -768 933 -672
rect 987 -701 993 -341
rect 772 -817 912 -813
rect 917 -817 932 -813
rect 772 -822 777 -817
rect 650 -823 777 -822
rect 527 -827 777 -823
rect 527 -832 532 -827
rect 402 -836 532 -832
rect 408 -849 412 -836
rect 424 -849 428 -836
rect 462 -849 466 -836
rect 482 -849 486 -836
rect 570 -840 574 -827
rect 586 -840 590 -827
rect 624 -840 628 -827
rect 644 -840 648 -827
rect 807 -830 811 -817
rect 823 -830 827 -817
rect 861 -830 865 -817
rect 881 -830 885 -817
rect 416 -874 420 -855
rect 443 -865 447 -855
rect 394 -878 409 -874
rect 416 -878 435 -874
rect 270 -886 402 -882
rect 270 -888 276 -886
rect 416 -897 420 -878
rect 443 -897 447 -870
rect 474 -874 478 -855
rect 578 -865 582 -846
rect 605 -856 609 -846
rect 516 -866 571 -865
rect 509 -869 571 -866
rect 578 -869 597 -865
rect 509 -870 545 -869
rect 465 -878 478 -874
rect 474 -897 478 -878
rect 485 -881 489 -874
rect 516 -879 522 -873
rect 485 -893 489 -886
rect 408 -915 412 -901
rect 424 -915 428 -901
rect 462 -915 466 -901
rect 482 -915 486 -901
rect 403 -919 489 -915
rect 516 -921 521 -915
rect 539 -970 545 -870
rect 557 -877 564 -873
rect 557 -878 561 -877
rect 578 -888 582 -869
rect 605 -888 609 -861
rect 636 -865 640 -846
rect 676 -857 784 -855
rect 671 -859 784 -857
rect 815 -855 819 -836
rect 842 -846 846 -836
rect 789 -859 808 -855
rect 815 -859 834 -855
rect 671 -861 680 -859
rect 627 -869 640 -865
rect 636 -888 640 -869
rect 647 -872 651 -865
rect 647 -884 651 -877
rect 777 -867 801 -863
rect 570 -906 574 -892
rect 586 -906 590 -892
rect 624 -906 628 -892
rect 644 -906 648 -892
rect 656 -906 661 -904
rect 565 -910 661 -906
rect 777 -916 781 -867
rect 815 -878 819 -859
rect 842 -878 846 -851
rect 873 -855 877 -836
rect 954 -851 960 -846
rect 864 -859 877 -855
rect 873 -878 877 -859
rect 884 -862 888 -855
rect 884 -874 888 -867
rect 807 -896 811 -882
rect 823 -896 827 -882
rect 861 -896 865 -882
rect 881 -896 885 -882
rect 807 -900 892 -896
rect 570 -920 781 -916
rect 690 -941 754 -938
rect 696 -956 700 -941
rect 715 -956 719 -941
rect 739 -956 743 -941
rect 705 -970 709 -962
rect 747 -970 751 -962
rect 777 -969 781 -920
rect 821 -940 909 -937
rect 824 -955 828 -940
rect 843 -955 847 -940
rect 867 -955 871 -940
rect 917 -940 932 -937
rect 833 -969 837 -961
rect 875 -969 879 -961
rect 757 -970 770 -969
rect 539 -974 697 -970
rect 705 -974 740 -970
rect 747 -974 770 -970
rect 777 -973 825 -969
rect 833 -973 868 -969
rect 875 -973 932 -969
rect 540 -975 689 -974
rect 669 -983 707 -979
rect 715 -988 719 -974
rect 747 -988 751 -974
rect 667 -999 691 -998
rect 696 -999 700 -992
rect 739 -999 743 -992
rect 667 -1002 753 -999
rect 763 -1049 770 -974
rect 789 -982 835 -978
rect 843 -987 847 -973
rect 875 -987 879 -973
rect 824 -998 828 -991
rect 867 -998 871 -991
rect 821 -1001 886 -998
rect 859 -1015 909 -1010
rect 865 -1027 869 -1015
rect 893 -1027 897 -1015
rect 819 -1046 866 -1042
rect 819 -1090 823 -1046
rect 883 -1047 887 -1033
rect 901 -1047 905 -1033
rect 862 -1053 876 -1049
rect 883 -1051 894 -1047
rect 901 -1051 917 -1047
rect 883 -1057 887 -1051
rect 874 -1061 887 -1057
rect 874 -1065 878 -1061
rect 901 -1065 905 -1051
rect 865 -1076 869 -1069
rect 883 -1076 887 -1069
rect 893 -1076 897 -1069
rect 861 -1081 907 -1076
rect 928 -1090 932 -973
rect 956 -1051 961 -1046
rect 987 -1076 993 -707
rect 1032 -429 1040 -63
rect 1032 -796 1040 -434
rect 819 -1095 932 -1090
<< m2contact >>
rect 385 202 390 207
rect 344 186 349 191
rect 547 211 552 216
rect 446 202 451 207
rect 464 193 471 199
rect 426 186 431 191
rect 493 193 499 199
rect 506 195 511 200
rect 608 211 613 216
rect 726 213 731 218
rect 784 221 789 226
rect 588 195 593 200
rect 743 205 748 210
rect 891 221 896 226
rect 825 205 830 210
rect 603 87 611 94
rect 726 90 731 95
rect 705 17 713 23
rect 797 17 804 23
rect 859 21 864 26
rect 852 -9 859 -4
rect 893 21 898 26
rect 868 -77 873 -72
rect 394 -130 399 -125
rect 353 -146 358 -141
rect 556 -121 561 -116
rect 455 -130 460 -125
rect 473 -139 480 -133
rect 435 -146 440 -141
rect 502 -139 508 -133
rect 515 -137 520 -132
rect 617 -121 622 -116
rect 735 -119 740 -114
rect 793 -111 798 -106
rect 597 -137 602 -132
rect 752 -127 757 -122
rect 900 -111 905 -106
rect 834 -127 839 -122
rect 612 -245 620 -238
rect 735 -242 740 -237
rect 714 -315 722 -309
rect 806 -315 813 -309
rect 868 -311 873 -306
rect 902 -311 907 -306
rect 1032 -63 1040 -58
rect 884 -434 889 -429
rect 415 -496 420 -491
rect 374 -512 379 -507
rect 577 -487 582 -482
rect 476 -496 481 -491
rect 494 -505 501 -499
rect 456 -512 461 -507
rect 523 -505 529 -499
rect 536 -503 541 -498
rect 638 -487 643 -482
rect 756 -485 761 -480
rect 814 -477 819 -472
rect 618 -503 623 -498
rect 773 -493 778 -488
rect 921 -477 926 -472
rect 855 -493 860 -488
rect 633 -611 641 -604
rect 756 -608 761 -603
rect 735 -681 743 -675
rect 827 -681 834 -675
rect 889 -677 894 -672
rect 923 -677 928 -672
rect 912 -817 917 -811
rect 443 -870 448 -865
rect 402 -886 407 -881
rect 605 -861 610 -856
rect 504 -870 509 -865
rect 522 -879 529 -873
rect 484 -886 489 -881
rect 551 -879 557 -873
rect 564 -877 569 -872
rect 666 -861 671 -856
rect 784 -859 789 -854
rect 842 -851 847 -846
rect 646 -877 651 -872
rect 801 -867 806 -862
rect 949 -851 954 -846
rect 883 -867 888 -862
rect 661 -985 669 -978
rect 784 -982 789 -977
rect 763 -1055 771 -1049
rect 855 -1055 862 -1049
rect 917 -1051 922 -1046
rect 907 -1081 915 -1076
rect 951 -1051 956 -1046
rect 1032 -434 1040 -429
rect 1032 -801 1040 -796
rect 987 -1081 994 -1076
<< metal2 >>
rect 789 221 891 225
rect 552 211 608 215
rect 390 202 446 206
rect 471 193 493 199
rect 511 195 588 200
rect 349 186 426 191
rect 493 94 499 193
rect 726 95 731 213
rect 748 205 825 210
rect 493 87 603 94
rect 726 89 731 90
rect 713 17 797 23
rect 864 21 893 25
rect 859 -9 987 -4
rect 868 -63 1032 -60
rect 868 -72 873 -63
rect 798 -111 900 -107
rect 561 -121 617 -117
rect 399 -130 455 -126
rect 480 -139 502 -133
rect 520 -137 597 -132
rect 358 -146 435 -141
rect 502 -238 508 -139
rect 735 -237 740 -119
rect 757 -127 834 -122
rect 502 -245 612 -238
rect 735 -243 740 -242
rect 722 -315 806 -309
rect 873 -311 902 -307
rect 860 -341 987 -336
rect 889 -434 1032 -429
rect 819 -477 921 -473
rect 582 -487 638 -483
rect 420 -496 476 -492
rect 501 -505 523 -499
rect 541 -503 618 -498
rect 379 -512 456 -507
rect 523 -604 529 -505
rect 756 -603 761 -485
rect 778 -493 855 -488
rect 523 -611 633 -604
rect 756 -609 761 -608
rect 743 -681 827 -675
rect 894 -677 923 -673
rect 880 -707 987 -702
rect 912 -801 1032 -797
rect 912 -811 917 -801
rect 847 -851 949 -847
rect 610 -861 666 -857
rect 448 -870 504 -866
rect 529 -879 551 -873
rect 569 -877 646 -872
rect 407 -886 484 -881
rect 551 -978 557 -879
rect 784 -977 789 -859
rect 806 -867 883 -862
rect 551 -985 661 -978
rect 784 -983 789 -982
rect 771 -1055 855 -1049
rect 922 -1051 951 -1047
rect 915 -1081 987 -1076
<< m123contact >>
rect 874 254 880 259
rect 430 152 436 157
rect 463 151 471 157
rect 603 162 608 168
rect 507 151 512 157
rect 696 131 701 136
rect 744 171 749 177
rect 755 131 763 136
rect 851 131 859 136
rect 874 132 882 137
rect 603 70 608 75
rect 695 70 700 75
rect 758 70 763 75
rect 851 56 859 62
rect 793 -9 803 -4
rect 987 -9 994 -4
rect 898 -37 903 -32
rect 883 -78 889 -73
rect 442 -179 447 -174
rect 472 -181 480 -175
rect 612 -170 617 -164
rect 516 -181 521 -175
rect 705 -201 710 -196
rect 753 -160 758 -155
rect 764 -201 772 -196
rect 860 -201 868 -196
rect 883 -200 890 -195
rect 612 -262 617 -257
rect 704 -262 709 -257
rect 767 -262 772 -257
rect 860 -276 868 -270
rect 802 -341 812 -336
rect 987 -341 995 -336
rect 905 -406 912 -398
rect 904 -444 910 -439
rect 461 -546 467 -540
rect 493 -547 501 -541
rect 633 -536 638 -530
rect 537 -547 542 -541
rect 726 -567 731 -562
rect 774 -526 779 -521
rect 785 -567 793 -562
rect 881 -567 889 -562
rect 904 -566 911 -561
rect 633 -628 638 -622
rect 725 -628 730 -623
rect 788 -628 793 -623
rect 881 -642 889 -636
rect 823 -707 833 -702
rect 987 -707 993 -701
rect 927 -774 933 -768
rect 932 -819 938 -813
rect 489 -920 494 -915
rect 521 -921 529 -915
rect 661 -910 666 -904
rect 565 -921 570 -915
rect 754 -941 759 -936
rect 802 -900 807 -895
rect 813 -941 821 -936
rect 909 -941 917 -936
rect 932 -940 939 -934
rect 661 -1002 667 -997
rect 753 -1002 759 -997
rect 816 -1002 821 -997
rect 909 -1016 917 -1010
rect 851 -1081 861 -1076
<< metal3 >>
rect 744 167 749 171
rect 608 163 749 167
rect 430 75 436 152
rect 471 151 507 157
rect 603 75 608 162
rect 874 137 880 254
rect 701 131 755 135
rect 430 70 603 75
rect 700 70 758 73
rect 731 -4 735 70
rect 851 62 858 131
rect 731 -9 793 -4
rect 479 -37 898 -32
rect 480 -175 486 -37
rect 753 -165 758 -160
rect 617 -169 758 -165
rect 442 -257 447 -179
rect 480 -181 516 -175
rect 612 -257 617 -170
rect 883 -195 889 -78
rect 710 -201 764 -197
rect 442 -262 612 -257
rect 709 -262 767 -259
rect 442 -264 447 -262
rect 740 -336 744 -262
rect 860 -270 867 -201
rect 740 -341 802 -336
rect 501 -406 905 -398
rect 502 -541 508 -406
rect 774 -531 779 -526
rect 638 -535 779 -531
rect 461 -623 467 -546
rect 501 -547 537 -541
rect 633 -622 638 -536
rect 904 -561 910 -444
rect 731 -567 785 -563
rect 461 -628 633 -623
rect 730 -628 788 -625
rect 761 -702 765 -628
rect 881 -636 888 -567
rect 761 -707 823 -702
rect 539 -774 927 -768
rect 539 -915 546 -774
rect 802 -905 807 -900
rect 666 -909 807 -905
rect 489 -997 494 -920
rect 529 -921 565 -915
rect 661 -997 666 -910
rect 932 -934 938 -819
rect 759 -941 813 -937
rect 489 -1002 661 -997
rect 759 -1002 816 -999
rect 789 -1076 793 -1002
rect 909 -1010 916 -941
rect 789 -1081 851 -1076
<< labels >>
rlabel metal1 336 186 342 190 3 B0
rlabel metal1 458 193 464 199 1 A0
rlabel metal1 458 151 463 157 1 M
rlabel metal1 896 221 902 226 1 S0
rlabel metal1 467 -139 473 -133 1 A1
rlabel metal1 345 -146 350 -142 1 B1
rlabel metal1 905 -111 911 -106 1 S1
rlabel metal1 488 -505 494 -499 1 A2
rlabel metal1 366 -512 370 -508 1 B2
rlabel metal1 394 -878 399 -874 1 B3
rlabel metal1 516 -879 522 -873 1 A3
rlabel metal1 954 -851 960 -846 7 S3
rlabel metal1 926 -477 932 -472 1 S2
rlabel metal1 956 -1051 961 -1046 7 Carryout
rlabel metal1 336 194 342 198 3 M
rlabel metal1 345 -138 350 -134 1 M
rlabel metal1 366 -504 370 -500 1 M
rlabel metal1 394 -886 399 -882 1 M
rlabel metal1 907 -311 912 -306 1 Carry1
rlabel metal1 928 -677 933 -672 1 Carry2
rlabel metal1 672 -119 686 -115 1 D1
rlabel metal1 467 -181 472 -175 1 Carry0
rlabel metal1 516 -921 521 -915 1 Carry2
rlabel metal1 344 236 434 240 1 VDD
rlabel metal1 506 245 536 249 1 VDD
rlabel metal1 743 255 833 259 5 VDD
rlabel metal1 533 -87 547 -83 1 VDD
rlabel metal1 777 -77 791 -73 1 VDD
rlabel metal1 804 -200 811 -197 1 VDD
rlabel metal1 374 -462 464 -458 1 VDD
rlabel metal1 773 -443 863 -439 5 VDD
rlabel metal1 536 -453 566 -449 1 VDD
rlabel metal1 402 -836 492 -832 1 VDD
rlabel metal1 564 -827 594 -823 1 VDD
rlabel metal1 801 -817 891 -813 5 VDD
rlabel metal1 507 162 597 166 1 GND
rlabel metal1 522 -170 536 -166 1 GND
rlabel metal1 783 -160 797 -156 1 GND
rlabel metal1 799 -261 806 -258 1 GND
rlabel metal1 537 -536 627 -532 1 GND
rlabel metal1 379 154 381 157 1 GND
rlabel metal1 376 -95 382 -92 1 VDD
rlabel metal1 383 -179 389 -176 1 GND
rlabel metal1 614 -909 621 -906 1 GND
rlabel metal1 838 -900 845 -897 1 GND
rlabel metal1 1032 132 1040 146 7 VDD
rlabel metal1 987 -275 993 -267 1 GND
rlabel metal1 769 173 776 176 1 GND
<< end >>
