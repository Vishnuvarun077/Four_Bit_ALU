magic
tech scmos
timestamp 1701449652
<< nwell >>
rect 601 32 638 50
rect 644 32 668 50
rect 687 32 724 50
rect 730 32 754 50
rect 777 32 814 50
rect 820 32 844 50
rect 872 32 909 50
rect 915 32 939 50
rect 956 32 993 50
rect 999 32 1023 50
rect 1042 32 1079 50
rect 1085 32 1109 50
rect 1132 32 1169 50
rect 1175 32 1199 50
rect 1227 32 1264 50
rect 1270 32 1294 50
<< ntransistor >>
rect 612 8 614 12
rect 622 8 624 12
rect 655 8 657 12
rect 698 8 700 12
rect 708 8 710 12
rect 741 8 743 12
rect 788 8 790 12
rect 798 8 800 12
rect 831 8 833 12
rect 883 8 885 12
rect 893 8 895 12
rect 926 8 928 12
rect 967 8 969 12
rect 977 8 979 12
rect 1010 8 1012 12
rect 1053 8 1055 12
rect 1063 8 1065 12
rect 1096 8 1098 12
rect 1143 8 1145 12
rect 1153 8 1155 12
rect 1186 8 1188 12
rect 1238 8 1240 12
rect 1248 8 1250 12
rect 1281 8 1283 12
<< ptransistor >>
rect 612 38 614 44
rect 622 38 624 44
rect 655 38 657 44
rect 698 38 700 44
rect 708 38 710 44
rect 741 38 743 44
rect 788 38 790 44
rect 798 38 800 44
rect 831 38 833 44
rect 883 38 885 44
rect 893 38 895 44
rect 926 38 928 44
rect 967 38 969 44
rect 977 38 979 44
rect 1010 38 1012 44
rect 1053 38 1055 44
rect 1063 38 1065 44
rect 1096 38 1098 44
rect 1143 38 1145 44
rect 1153 38 1155 44
rect 1186 38 1188 44
rect 1238 38 1240 44
rect 1248 38 1250 44
rect 1281 38 1283 44
<< ndiffusion >>
rect 611 8 612 12
rect 614 8 622 12
rect 624 8 626 12
rect 654 8 655 12
rect 657 8 658 12
rect 697 8 698 12
rect 700 8 708 12
rect 710 8 712 12
rect 740 8 741 12
rect 743 8 744 12
rect 787 8 788 12
rect 790 8 798 12
rect 800 8 802 12
rect 830 8 831 12
rect 833 8 834 12
rect 882 8 883 12
rect 885 8 893 12
rect 895 8 897 12
rect 925 8 926 12
rect 928 8 929 12
rect 966 8 967 12
rect 969 8 977 12
rect 979 8 981 12
rect 1009 8 1010 12
rect 1012 8 1013 12
rect 1052 8 1053 12
rect 1055 8 1063 12
rect 1065 8 1067 12
rect 1095 8 1096 12
rect 1098 8 1099 12
rect 1142 8 1143 12
rect 1145 8 1153 12
rect 1155 8 1157 12
rect 1185 8 1186 12
rect 1188 8 1189 12
rect 1237 8 1238 12
rect 1240 8 1248 12
rect 1250 8 1252 12
rect 1280 8 1281 12
rect 1283 8 1284 12
<< pdiffusion >>
rect 611 38 612 44
rect 614 38 616 44
rect 620 38 622 44
rect 624 38 626 44
rect 654 38 655 44
rect 657 38 658 44
rect 697 38 698 44
rect 700 38 702 44
rect 706 38 708 44
rect 710 38 712 44
rect 740 38 741 44
rect 743 38 744 44
rect 787 38 788 44
rect 790 38 792 44
rect 796 38 798 44
rect 800 38 802 44
rect 830 38 831 44
rect 833 38 834 44
rect 882 38 883 44
rect 885 38 887 44
rect 891 38 893 44
rect 895 38 897 44
rect 925 38 926 44
rect 928 38 929 44
rect 966 38 967 44
rect 969 38 971 44
rect 975 38 977 44
rect 979 38 981 44
rect 1009 38 1010 44
rect 1012 38 1013 44
rect 1052 38 1053 44
rect 1055 38 1057 44
rect 1061 38 1063 44
rect 1065 38 1067 44
rect 1095 38 1096 44
rect 1098 38 1099 44
rect 1142 38 1143 44
rect 1145 38 1147 44
rect 1151 38 1153 44
rect 1155 38 1157 44
rect 1185 38 1186 44
rect 1188 38 1189 44
rect 1237 38 1238 44
rect 1240 38 1242 44
rect 1246 38 1248 44
rect 1250 38 1252 44
rect 1280 38 1281 44
rect 1283 38 1284 44
<< ndcontact >>
rect 607 8 611 12
rect 626 8 630 12
rect 650 8 654 12
rect 658 8 662 12
rect 693 8 697 12
rect 712 8 716 12
rect 736 8 740 12
rect 744 8 748 12
rect 783 8 787 12
rect 802 8 806 12
rect 826 8 830 12
rect 834 8 838 12
rect 878 8 882 12
rect 897 8 901 12
rect 921 8 925 12
rect 929 8 933 12
rect 962 8 966 12
rect 981 8 985 12
rect 1005 8 1009 12
rect 1013 8 1017 12
rect 1048 8 1052 12
rect 1067 8 1071 12
rect 1091 8 1095 12
rect 1099 8 1103 12
rect 1138 8 1142 12
rect 1157 8 1161 12
rect 1181 8 1185 12
rect 1189 8 1193 12
rect 1233 8 1237 12
rect 1252 8 1256 12
rect 1276 8 1280 12
rect 1284 8 1288 12
<< pdcontact >>
rect 607 38 611 44
rect 616 38 620 44
rect 626 38 630 44
rect 650 38 654 44
rect 658 38 662 44
rect 693 38 697 44
rect 702 38 706 44
rect 712 38 716 44
rect 736 38 740 44
rect 744 38 748 44
rect 783 38 787 44
rect 792 38 796 44
rect 802 38 806 44
rect 826 38 830 44
rect 834 38 838 44
rect 878 38 882 44
rect 887 38 891 44
rect 897 38 901 44
rect 921 38 925 44
rect 929 38 933 44
rect 962 38 966 44
rect 971 38 975 44
rect 981 38 985 44
rect 1005 38 1009 44
rect 1013 38 1017 44
rect 1048 38 1052 44
rect 1057 38 1061 44
rect 1067 38 1071 44
rect 1091 38 1095 44
rect 1099 38 1103 44
rect 1138 38 1142 44
rect 1147 38 1151 44
rect 1157 38 1161 44
rect 1181 38 1185 44
rect 1189 38 1193 44
rect 1233 38 1237 44
rect 1242 38 1246 44
rect 1252 38 1256 44
rect 1276 38 1280 44
rect 1284 38 1288 44
<< polysilicon >>
rect 612 44 614 53
rect 622 44 624 53
rect 655 44 657 53
rect 698 44 700 53
rect 708 44 710 53
rect 741 44 743 53
rect 788 44 790 53
rect 798 44 800 53
rect 831 44 833 53
rect 883 44 885 53
rect 893 44 895 53
rect 926 44 928 53
rect 967 44 969 53
rect 977 44 979 53
rect 1010 44 1012 53
rect 1053 44 1055 53
rect 1063 44 1065 53
rect 1096 44 1098 53
rect 1143 44 1145 53
rect 1153 44 1155 53
rect 1186 44 1188 53
rect 1238 44 1240 53
rect 1248 44 1250 53
rect 1281 44 1283 53
rect 612 12 614 38
rect 622 12 624 38
rect 655 12 657 38
rect 698 12 700 38
rect 708 12 710 38
rect 741 12 743 38
rect 788 12 790 38
rect 798 12 800 38
rect 831 12 833 38
rect 883 12 885 38
rect 893 12 895 38
rect 926 12 928 38
rect 967 12 969 38
rect 977 12 979 38
rect 1010 12 1012 38
rect 1053 12 1055 38
rect 1063 12 1065 38
rect 1096 12 1098 38
rect 1143 12 1145 38
rect 1153 12 1155 38
rect 1186 12 1188 38
rect 1238 12 1240 38
rect 1248 12 1250 38
rect 1281 12 1283 38
rect 612 5 614 8
rect 622 5 624 8
rect 655 5 657 8
rect 698 5 700 8
rect 708 5 710 8
rect 741 5 743 8
rect 788 5 790 8
rect 798 5 800 8
rect 831 5 833 8
rect 883 5 885 8
rect 893 5 895 8
rect 926 5 928 8
rect 967 5 969 8
rect 977 5 979 8
rect 1010 5 1012 8
rect 1053 5 1055 8
rect 1063 5 1065 8
rect 1096 5 1098 8
rect 1143 5 1145 8
rect 1153 5 1155 8
rect 1186 5 1188 8
rect 1238 5 1240 8
rect 1248 5 1250 8
rect 1281 5 1283 8
<< polycontact >>
rect 608 26 612 30
rect 618 17 622 21
rect 651 26 655 30
rect 694 26 698 30
rect 704 17 708 21
rect 737 26 741 30
rect 784 26 788 30
rect 794 17 798 21
rect 827 26 831 30
rect 879 26 883 30
rect 889 17 893 21
rect 922 26 926 30
rect 963 26 967 30
rect 973 17 977 21
rect 1006 26 1010 30
rect 1049 26 1053 30
rect 1059 17 1063 21
rect 1092 26 1096 30
rect 1139 26 1143 30
rect 1149 17 1153 21
rect 1182 26 1186 30
rect 1234 26 1238 30
rect 1244 17 1248 21
rect 1277 26 1281 30
<< metal1 >>
rect 584 70 590 75
rect 601 59 1294 62
rect 607 44 611 59
rect 626 44 630 59
rect 650 44 654 59
rect 693 44 697 59
rect 712 44 716 59
rect 736 44 740 59
rect 783 44 787 59
rect 802 44 806 59
rect 826 44 830 59
rect 878 44 882 59
rect 897 44 901 59
rect 921 44 925 59
rect 962 44 966 59
rect 981 44 985 59
rect 1005 44 1009 59
rect 1048 44 1052 59
rect 1067 44 1071 59
rect 1091 44 1095 59
rect 1138 44 1142 59
rect 1157 44 1161 59
rect 1181 44 1185 59
rect 1233 44 1237 59
rect 1252 44 1256 59
rect 1276 44 1280 59
rect 616 30 620 38
rect 658 30 662 38
rect 702 30 706 38
rect 744 30 748 38
rect 792 30 796 38
rect 834 30 838 38
rect 887 30 891 38
rect 929 30 933 38
rect 971 30 975 38
rect 1013 30 1017 38
rect 1057 30 1061 38
rect 1099 30 1103 38
rect 1147 30 1151 38
rect 1189 30 1193 38
rect 1242 30 1246 38
rect 1284 30 1288 38
rect 596 26 608 30
rect 616 26 651 30
rect 658 26 671 30
rect 682 26 694 30
rect 702 26 737 30
rect 744 26 757 30
rect 772 26 784 30
rect 792 26 827 30
rect 834 26 847 30
rect 867 26 879 30
rect 887 26 922 30
rect 929 26 942 30
rect 951 26 963 30
rect 971 26 1006 30
rect 1013 26 1026 30
rect 1037 26 1049 30
rect 1057 26 1092 30
rect 1099 26 1112 30
rect 1127 26 1139 30
rect 1147 26 1182 30
rect 1189 26 1202 30
rect 1222 26 1234 30
rect 1242 26 1277 30
rect 1284 26 1297 30
rect 596 17 618 21
rect 626 12 630 26
rect 658 12 662 26
rect 681 17 704 21
rect 712 12 716 26
rect 744 12 748 26
rect 771 17 794 21
rect 802 12 806 26
rect 834 12 838 26
rect 865 17 889 21
rect 897 12 901 26
rect 929 12 933 26
rect 951 17 973 21
rect 981 12 985 26
rect 1013 12 1017 26
rect 1036 17 1059 21
rect 1067 12 1071 26
rect 1099 12 1103 26
rect 1126 17 1149 21
rect 1157 12 1161 26
rect 1189 12 1193 26
rect 1220 17 1244 21
rect 1252 12 1256 26
rect 1284 12 1288 26
rect 607 1 611 8
rect 650 1 654 8
rect 693 1 697 8
rect 736 1 740 8
rect 783 1 787 8
rect 826 1 830 8
rect 878 1 882 8
rect 921 1 925 8
rect 962 1 966 8
rect 1005 1 1009 8
rect 1048 1 1052 8
rect 1091 1 1095 8
rect 1138 1 1142 8
rect 1181 1 1185 8
rect 1233 1 1237 8
rect 1276 1 1280 8
rect 600 -2 1295 1
<< m2contact >>
rect 590 70 596 75
rect 590 16 596 21
rect 675 17 681 22
rect 765 17 771 22
rect 860 16 865 21
rect 945 16 951 21
rect 1030 17 1036 22
rect 1120 17 1126 22
rect 1215 16 1220 21
<< metal2 >>
rect 596 70 1220 75
rect 590 21 596 70
rect 675 22 681 70
rect 765 22 771 70
rect 860 21 865 70
rect 945 21 951 70
rect 1030 22 1036 70
rect 1120 22 1126 70
rect 1215 21 1220 70
<< labels >>
rlabel metal1 596 26 600 30 3 A0
rlabel metal1 682 26 686 30 1 A1
rlabel metal1 772 26 776 30 1 A2
rlabel metal1 867 26 871 30 1 A3
rlabel metal1 584 70 590 75 4 E
rlabel metal1 1229 -2 1239 1 1 GND
rlabel metal1 1241 59 1251 62 5 VDD
rlabel metal1 951 26 955 30 1 B0
rlabel metal1 1037 26 1041 30 1 B1
rlabel metal1 1127 26 1131 30 1 B2
rlabel metal1 1222 26 1226 30 1 B3
<< end >>
